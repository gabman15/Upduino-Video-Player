library IEEE;
use IEEE.STD_LOGIC_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.all;

entity scale_clock is
  port (
    clk_12Mhz : in  std_logic;
    rst       : in  std_logic;
    clk_10Hz   : out std_logic);
end scale_clock;

architecture Behavioral of scale_clock is

  signal prescaler : unsigned(23 downto 0);
  signal clk_10Hz_i : std_logic;
begin

  gen_clk : process (clk_12Mhz, rst)
  begin  -- process gen_clk
    if rst = '1' then
      clk_10Hz_i   <= '0';
      prescaler   <= (others => '0');
    elsif rising_edge(clk_12Mhz) then   -- rising clock edge
      if prescaler = X"124F80" then     -- 1 200 000 in hex
        prescaler   <= (others => '0');
        clk_10Hz_i   <= not clk_10Hz_i;
      else
        prescaler <= prescaler + "1";
      end if;
    end if;
  end process gen_clk;

clk_10Hz <= clk_10Hz_i;

end Behavioral;
