library IEEE;
use IEEE.std_logic_1164.all;
entity rom is
port(
clk : in std_logic;
addr : in std_logic_vector (10 downto 0);
data : out std_logic_vector (767 downto 0)
);
end rom;
architecture synth of rom is
begin
process(clk) is
begin
if rising_edge(clk) then
case addr is
 when "00000000000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000100" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000000111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001100" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000010000" => data <= 768x"000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000001000000030000000100000003000000030000000300000001000000000000000000000000000000000000000000000000";
 when "00000010001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000080000000c00000008000000050000000f000000170000001f0000001f0000000f00000007000000030000000300000003000000010000000100000001";
 when "00000010010" => data <= 768x"0000003f0000005f0000003f0000001f0000003f0000001f0000001f0000001f0000003f0000001f0000003f0000007f0000003f0000005f0000003f0000007f0000003f0000005f0000003f0000001f0000003f0000001f0000000f00000017";
 when "00000010011" => data <= 768x"00000fff00000fff00000fff000007ff00000fff00000fff00000fff000017ff00000fff000007ff00000fff0000077f00000fff000007ff000007ff000001ff000001ff000000ff000000ff0000007f0000007f0000007f0000003f0000001f";
 when "00000010100" => data <= 768x"000003ff000005ff000003ff0000077f00000fff00001fff00001fff000015ff000003ff000001ff000003ff0000017f0000007f0000001f0000001f0000001f0000001f0000001f0000000f0000001f0000000f000000070000000300000011";
 when "00000010101" => data <= 768x"000000ff000001ff000001ff0000017f000003ff000007ff000003ff4000007f400000ffc000007f8000003f0000001f0000000f0000000700000007000000070000000700000007000000070000000700000003000000010000000000000000";
 when "00000010110" => data <= 768x"f000007ff000007ff000007ff000007fe000007ff000007fe00000fff010017fe020007fd000007fe000003fc000001fe000000fc0000007c0000007c00000078000000700000007000000070000000700000003000000000000000000000000";
 when "00000010111" => data <= 768x"f800000ffc00005ffe00003fff00003ffe00003ffc40007ffe00003ff400007ffe00003ffc04007ffe00007ffc00007ffe00003ffc00001ff800000ff0000007f0000007f0000007e0000007c0000007c0000003c00000008000000010000000";
 when "00000011000" => data <= 768x"ff00000fff00001fff80003f7f00001fff80003fff00001fff80003fff100017ff80003fff00001fff80003f7f00001fff80000fff000007ff000007ff000007fe000007fc000007f800000370000001f8000000f0000000e0000000f0000001";
 when "00000011001" => data <= 768x"ff80001fffc0001fffe0003f7f40001fffc0003fffc4001fffc8003fffc0001fffc8003fffd0005fffc0000f7fc00007ffc00007ffc00007ffc00007ffc00007ff000003ff000005fe0000007f000000fe000000fc000001fc000000fc000000";
 when "00000011010" => data <= 768x"fff0001ffff0001ffff0003f7f70001fffe0003ffff0007fffe0003fff700017ffe0003ffff4001ffff0000f7f700007ffe00003fff00007ffe00003ffc00007ff800003ffc00000ff8000007f000001ff800020ff000040ff000020ff000040";
 when "00000011011" => data <= 768x"fff0000ffff00007fff8001f7f70001ffff8003ffffc001ffff8003ffff00077fff8003ffff0001ffff8001f7f700017fff80007fff00007fff00007ffd00007ffc00007ffc00005ffe000017f400001ffc00003ffc00001ff800003ff000041";
 when "00000011100" => data <= 768x"ffe0003ffff0001ffff8003f7f71007ffff8003ffffc007ffffc003ffff4003ffffc003ffffc007ffff8007fff71001ffff0001ffff0001fffe0001fffc0001fffc0000fffc00007ffe000077fc00007ff80000fffc00007ff800007ff000007";
 when "00000011101" => data <= 768x"fff000fffff0007fffe000ff7f7001fffff800fffffc007ffff8007ffff4007ffff800fffff0007fffe000ffffc0007fffe0007fffc0007fff80007fff000017ff80001fffc0041fff80063f7f00041fff80061fff00041ffe00060fff000417";
 when "00000011110" => data <= 768x"ffe000ffffc001ffffc001ff7f70017ffff003fffff001fffff801fffff001f7fff001ffffd001ffffc001ff7fc001ffff8000ffffc0007fff80007fff00007fff80007fff00107fff00083f7f00117ffe00083ffe00107ffe00083ff4001017";
 when "00000011111" => data <= 768x"ffa000ffffc001ffffc003ff7fc0037fffe003fffff007ffffe007fffff007fffff003fffff007ffffc003ffffc001ffff8001ffffc001ffff8000fff700007fff00007fff00007ffe00007f7f00117ffe00007ffc00107ffc00007ff000107f";
 when "00000100000" => data <= 768x"ff8001ffffc001ffffe003ff7fc0077fffc007ffffc007ffffe00fffff5007ffffe00ffffff007ffffe00fffffc007ffff8003ffffc001ffff8001fff70001f7ff0001ffff0005fffe0000fffc00007ffc0020fffc00007ff80000fff000007f";
 when "00000100001" => data <= 768x"ff8003ffffc007ffffc007ff7fc0077fffe00fffffc01fffffc00fffffc01fffffe01fffffc01fffffc00fff7f0017ffff800fffff0007fffe0003fff70003f7fe0003fffc0001fffe0001fffc00017ffc0001fffc0001fff80000fff0000177";
 when "00000100010" => data <= 768x"ff0007ffff4007ffff800fff7f001f7fff801fffffc01fffffc01fffffc01fffffe03fffffc01fffff801fff7f001f7fff800fffff0007fffe000ffff70007f7fe2003fffc4007fffe2003ff7c00037ff80003fff84001fff80003fff00001ff";
 when "00000100011" => data <= 768x"ff000fffff401fffff800fff7f001f7fff803fffffc07fffffc03fffff4037ffffc03fffffc03fffff803fff7f001f7fff001fffff001ffffe000ffff70017f7fe200ffffc4007fffe2007ff7c00077ff80003fffc4007fff80003fff00001f7";
 when "00000100100" => data <= 768x"ff000fffff001fffff801fff7f001f7fff803fffffc07fffffc07fffffc077ffffc03fffffc07fffff803fff7f003f7fff803fffff001ffffe000ffff7001ff7ff000fffff0007fffe0007ff7c00077ffc0003fffc0007fff80003fffc0003f7";
 when "00000100101" => data <= 768x"ff800fffff0007ffff800fff7f401f7fffc03fffffc01fffffc03fffffc07fffffc07fffffc07fffffc01fff7fc01f7fff800fffff000fffff800fffff1007f7ff800fffff1007ffff0007ff7f10077ffe0003fffc0007fffe0003fffc0003f7";
 when "00000100110" => data <= 768x"ff8007ffffc007ffffc00fff7f701f7fffe01fffffc01fffffe03fffff407fffffe03fffffc01fffffc00fff7f40177fff800fffffc007ffff880fffffc007f7ff8807ffffc407ffff8803ff7f00017fff0003ffff1001ffff0003ffff1001ff";
 when "00000100111" => data <= 768x"ffc007ffffc007ffffe00fff7f701f7ffff00ffffff01ffffff01ffffff01fffffe03ffffff01fffffe00fff7fc0077fffc007ffffc007ffff8007ffff9007f7ff8003ffffc401ffff8001ff7fc401ffff8001ffffc401ffff8001ffffd001ff";
 when "00000101000" => data <= 768x"fffb07ffffc007ffffe007ff7f70177ffff00ffffff007fffff80ffffff01ffffff01ffffff01ffffff00fff7f70077fffe007ffffc007ffffc003ffffd003f7ffb003ffffd001ffff8000ff7f40017fffa000ffffc001ffffe000ffffc001ff";
 when "00000101001" => data <= 768x"fffb87ffffd007ffffe007ff7f70177ffff00ffffff007fffff80ffff7f017fffff80ffffffc0ffffff80fff7f70077fffe007ffffc007ffffe803ffffd001f7ffd001ffffd001ffffc000ff7fd0017fffe000ffffc0007fffe000fffff0017f";
 when "00000101010" => data <= 768x"fffb83fffff007ffffe007ff7f70077ffff807fffffc07fffffc0ffffffc17fffff80ffffffc07fffff807ff7f70077ffff003fffff401ffffe003ffff7011f7ffe001ffffc001ffffc000ff7fc0007fffe000fffff0007ffff000fffff0007f";
 when "00000101011" => data <= 768x"fff883fffff007fffff803ff7f71077ffffc07fffffc07fffffc0ffffffc07fffffc0ffffffc07fffffc03ff7f7c07fffff803fffff001fffff001fffff011f7fff001fffff001ffffe000ff7f70007fffe000fffff0007ffff800fffff0007f";
 when "00000101100" => data <= 768x"fffa83fffff001fffff803ff7f7c077ffffe03fffffc07fffffe0ffffff407fffffe07fffffc07fffffc03ff7f7c037ffff803fffffc01fffff803fffff011f7fff001fffff001ffffe000ff7ff0007fffe000fffff0007ffff800fffff0007f";
 when "00000101101" => data <= 768x"fffffbfffffd41fffff803ff7f70037ffff807fffffc07fffffe0ffff7ff07fffffe0ffffffc07fffffc07ff7f7c077ffff803fffffc01fffff803fffff011f7ffe001fffff001ffffe000ff7f60017fffe000fffff000fffff800fff7f0047f";
 when "00000101110" => data <= 768x"fffffffffff047fffff803ff7f70077ffff80ffffffc07fffffc0ffffff607fffffe0ffffffc07fffff807ff7f70077ffff803fffff017fffff003fffff01377ffe013ffffc011ffffe000ff7f4011ffffe001fffff001fffff008fffff005ff";
 when "00000101111" => data <= 768x"fffbfffffff047fffff807ff7f70077ffff80ffffffc1ffffffc0ffffffc17fffffc0ffffffc07fffff80fff7f70077ffff007fffff007ffffe027fffff03777ffe023ffffc011ffffc003ff7fc011ffffe003ffffc011ffffe009ffff6005ff";
 when "00000110000" => data <= 768x"fffbfffffff157fffff807ff7f71077ffff80ffffff41ffffff81ffffffc1ffffff81ffffff01ffffff80fff7f70077fffe007fffff047ffffe007ffffc047f7ffc027ffffc047ffffc003ff7fc0177fffc003ffffc017ffffc003ffffc013f7";
 when "00000110001" => data <= 768x"fffffffffff1dffffff00fff7f70077ffff80ffffff01ffffff81ffffff01ffffff83ffffff41ffffff81fff7f701f7fffe00ffffff007ffffe007ffffc057f7ffc007ffffc047ffff8007ff7f40077fff8003ffffc007ffffc007ffffc017f7";
 when "00000110010" => data <= 768x"fffffffffff1dffffff00fff7f70077ffff80ffffff01ffffff83ffffff03ffffff83ffffff01ffffff01fff7f701f7fffe00fffffc007ffffe00fffffc007f7ff8007ffffc007ffff8007ff7f00077fff8007ffffc007ffff800fffff8007f7";
 when "00000110011" => data <= 768x"fffffffffff15fffffe00fff7f701f7ffff01ffffff01ffffff83ffffff07ffffff03ffffff07fffffe03fff7f701f7fffe01fffffc01fffffc00fffffc017f7ff800fffff0007ffff800fff7f00077fff800fffff001fffff800fffff001ff7";
 when "00000110100" => data <= 768x"ffffffffffc55fffffe01fff7f701f7fffe03ffffff07ffffff03ffffff07ffffff03ffffff07fffffe03fff7f401f7fffe01fffffc01fffffc01fffffd01ff7ff800fffff000fffff800fff7f00177fff800fffff001fffff801fffff401ff7";
 when "00000110101" => data <= 768x"ffffffffffc55fffffe01fff7f401f7fffe03fffffc07fffffe07ffff7f07ffffff07ffffff07fffffe03fff7f403f7fffe03fffffc01fffffc01fffffd01ff7ff800fffff000fffff800fff7f001f7fff800fffff001fffff801fffff401ff7";
 when "00000110110" => data <= 768x"ffffffffffd55fffffe01fff7f401f7fffe03ffffff07fffffe07ffff7f07ffffff07ffffff07fffffe03fff7f701f7fffe03fffffc01fffffe01fffffc01ff7ff800fffff800fffff800fff7f001f7fff800fffff801fffffa00fffff401ff7";
 when "00000110111" => data <= 768x"fffffffffff55fffffe00fff7ff01f7ffff03ffffff01ffffff03fffff707ffffff03ffffff01fffffe01fff7ff01f7fffe01fffffe41fffffe40fffffc417f7ffc007ffffc407ffff880fff7fc0077fff800fffffd007ffff800ffffff007f7";
 when "00000111000" => data <= 768x"fffffffffff51fffffe00fff7f701f7ffff01ffffff01ffffff83ffffff07ffffff03ffffff01fffffe01fff7f701f7fffe00fffffc40fffffe00fffff5407f7ffe007ffffc407ffffc007ff7fc4077fffc807ffffd007ffffd007fffff007f7";
 when "00000111001" => data <= 768x"fffffffffff75fffffe00fff7f701f7ffff01ffffff01ffffff81ffffff017fffff83ffffff01ffffff00fff7f70177fffe00fffffd007ffffe007ffffd007f7ffe203ffffc401ffffe003ff7f4403ffffe003ffffc407ffffe807fffff007f7";
 when "00000111010" => data <= 768x"ffffffffffffdffffff80fff7f70177ffff00ffffffc1ffffff80ffffffc1ffffff81ffffffc1ffffff80fff7f7017fffff00ffffff007ffffe807fffff107ffffe003ffffc001ffffe003ff7f70017fffe003fffff401ffffe803fffff00777";
 when "00000111011" => data <= 768x"fffffffffffdc7fffff00fff7ff0077ffff80ffffffc07fffffc0ffffffc1ffffffc0ffffffc0ffffff80fff7ff1077ffff007fffff007ffffe003fffff003ffffe003ffffc001ffffe001ff7ff001fffff001fffff401fffff801fffff001ff";
 when "00000111100" => data <= 768x"fffffffffff547fffff807ff7f70077ffff80ffffffc07fffffc0ffffffc17fffffe0ffffffc07fffffc0fff7f7c077ffff803fffff017fffff003fffff011f7ffe001fffff001ffffe001ff7ff001fffff001fffff401fffff800fffff001ff";
 when "00000111101" => data <= 768x"ffffe7fffffd47fffff807ff7f7c07fffffc07fffffc07fffffe0ffffffc17fffffe0ffffffc07fffffc07ff7f7c077ffff803fffff007fffff003ffff7011f7ffe001fffff001ffffe001ff7f7001fffff001fffffc01fffff800fffff001f7";
 when "00000111110" => data <= 768x"fffffffffffdd7fffff803ff7f7c077ffffc07fffffc07fffffe0ffffff717fffffe0ffffffc07fffffe07ff7f7c077ffff803fffff007fffff003ffff7013f7ffe001ffffe001ffffe001ff7ff001fffff001fffff405fffff800fffff005f7";
 when "00000111111" => data <= 768x"fffffffffffd57fffff807ff7ff0077ffff80ffffffc07fffffe0fffffff07fffffe0ffffffc07fffffc0fff7f74077ffff803fffff017fffff003fffff013f7ffe003ffffc001ffffe001ff7f7001fffff001fffff005fffff004fffff005f7";
 when "00001000000" => data <= 768x"fffffffffff557fffff807ff7f7007fffff80ffffffc1ffffffc0ffffffc17fffffe0ffffffc1ffffff80fff7f70077ffff007fffff007ffffe027fffff007f7ffe023ffffc001ffffe003ff7f40117fffe003fffff001ffffe009fffff005f7";
 when "00001000001" => data <= 768x"fffffffffff157fffff807ff7f7007fffff80ffffffc1ffffffc1ffffffc1ffffff81ffffffc1ffffff80fff7f70077ffff007fffff047ffffe007ffffd047f7ffe023ffffc047ffffc003ff7fc0177fffe003ffffc017ffffe00bffffc007f7";
 when "00001000010" => data <= 768x"fffffffffff1fffffff00fff7f7007fffff80ffffff01ffffff81ffffff41ffffff81ffffffc1ffffff80fff7f701f7fffe00ffffff007ffffe007ffffc057f7ffc007ffffc047ffffc007ff7fc007ffffc007ffffc017ffffc007ffffc017f7";
 when "00001000011" => data <= 768x"fffffffffff5fffffff00fff7f7007fffff00ffffff01ffffff81ffffff01ffffff83ffffff01ffffff01fff7f701f7fffe00fffffe007ffffe00fffffc007f7ffc007ffffc047ffff8007ff7fc0077fff8007ffffc007ffff800fffffc017f7";
 when "00001000100" => data <= 768x"fffffffffff15ffffff007ff7f7007fffff80ffffff01ffffff81ffffff01ffffff81ffffff81ffffff81fff7f701f7ffff00ffffff007ffffe007fff7f007f7ffe003ffffc007ffff8003ff7f40037fff8003ffffc007ffff8007ffffc007f7";
 when "00001000101" => data <= 768x"fff3fffffff047fffff003ff7f70077ffff807fffff007fffff80ffffffc1ffffff80ffffffc1ffffff80fff7f70077ffff007fffff007ffffe003fff7f013ffffe003ffffc011ffffc001ff7fc011ffff8000ffffc001ffffc000ffffc001ff";
 when "00001000110" => data <= 768x"fff0fffffff041fffff001ff7f7001fffff803fffff005fffff803fffffc07fffff807fffffc07fffff807ff7f70077ffff803fffff005ffffe001fff7f001fffff000fffff0047fffe0087f7f70047fffe0003fffc0041fffc0003fffc0041f";
 when "00001000111" => data <= 768x"fffbfffffff050fffff000ff7f70007ffff800fffffc01fffff803fffffc01fffff803fffffc03fffff803ff7f7407fffff803fffff401fffff801fffff0017ffff0007ffff0007ffff8003f7f70041ffff8021ffff0071fffe0020fff70031f";
 when "00001001000" => data <= 768x"fffa383ffff0007ffff8003f7f7c003ffff8003ffffc007ffffc007ffffc007ffffc00fffffc01fffff800ff7f7d01fffffa01fffffc01fffffc00fffffc007ffffe003ffffc001ffffc000f7f740117fffe0307fffc0107fff80103fff00103";
 when "00001001001" => data <= 768x"ffff0a1ffffc001ffffe000f7f7f011ffffe000ffffc001ffffe001fffff0017ffff000fffff001ffffe803f7f7f007ffffe003fffff007ffffe007ff7f7007fffff003fffff0017fffe00077f770007fffe0003ffff0101fffe0081fffc0111";
 when "00001001010" => data <= 768x"fffffe1fffffc01fffff800f7f7f0007ffff000fffff000fffff000ff7f70007ffff8007ffffc007ffff800f7f7f9007ffff800fffffc00fffff800ff7ff801fffff803fffff001fffff000f7f7f0017ffff0003ffff0005ff9e0001f7000041";
 when "00001001011" => data <= 768x"fffffe3ffffff41fffffe03f7f7fc01fffff800fffff000fffff800fffff0007ffff8007ffffc007ffffc0077f7f4007ffffe007ffffc007ffffe007fff7c017ffffc00fffffc01fffff801f7f5f0017ff0f8007ff040007ff000007ff000007";
 when "00001001100" => data <= 768x"fffffffffffffc7ffffff8ff7f7f711fffffc01fffffc01fffff800fffff0017ffff800fffffc007ffffc0077f7f4007ffffe007fffff007ffffe007fff7f017ffffe00fffdfc05fff8f803f7f074037ff80002fffc0001fffe0000ffff00017";
 when "00001001101" => data <= 768x"fffffffffffff1fffffff8ff7f7f707fffffc03fffffc01fffff801fffff001fffff800fffffc01fffffc00f7f7f4007ffffe00ffffff007ffffe00ffffff017ffefe03fff07c05fff87c03f7f01003fff80002ffff0001ffff0001ffff0001f";
 when "00001001110" => data <= 768x"fffffffffffff1fffffff1ff7f7f717fffffc03fffffc01fffff801fffff001fffff800fffffc01fffffc00f7f7f401fffffe00ffffff01fffffe00fffd7f01fff8fe03fff07c07fff83803f7f41003fffe0003ffff0001fffe0001ffff0001f";
 when "00001001111" => data <= 768x"fffffffffffff7ffffffe3ff7f7f717fffffc03fffff801fffff803fffff001fffff001fffffc01fffffc01f7f7fc01fffffe01fffffe01fffffe01fffd7f01fff8fe03fff07c07fff80803f7fd0003fffe0001fffe0001fffe0003fffc0001f";
 when "00001010000" => data <= 768x"fffffffffffff7ffffffe3ff7f7f717fffff803fffff005fffff003fffff001fffff001fffff401fffff801f7f7fc01fffffe01fffffc01fffffe01fff57f05fff8f803fff05c07fff80803f7fd0007fffe0003fffc0001fffe0003fffc0001f";
 when "00001010001" => data <= 768x"ffffffffffffd7ffffffe7ff7f7fc07fffff807fffff007fffff003fffff0017ffff003fffff001fffff801f7f7fc01fffffe03fffffc01fffffe01fff57f05fff8f807fff05c07fff80807f7fd0007fffe0003fffc0001fffe0003fffc0001f";
 when "00001010010" => data <= 768x"ffffffffffffffffffffc7ff7f7f417fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff8f807fff05c07fff80807f7fd0007fffe0003fffc0005fffe0003fffc0001f";
 when "00001010011" => data <= 768x"ffffffffffffffffffffc7ff7f7f417fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff8f807fff07c07fff80807f7fd0007fffe0003ffff0005fffe0003fffe00017";
 when "00001010100" => data <= 768x"ffffffffffffd7ffffffc7ff7f7fc07fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff87a07fff05c07fff80807f7fd0007fffe0003ffff0005fffe0003ffff00017";
 when "00001010101" => data <= 768x"ffffffffffffd7ffffffc3ff7f7fc07fffff807fffff007fffff003fffff0017ffff003fffff001fffff801f7f7fc01fffffc01fffffc01fffffe03fff47e07fff87e07fffc5c07fff80807f7fd0007fffe0003ffff0005fffe0003ffff00017";
 when "00001010110" => data <= 768x"ffffffffffffc7ffffffc2ff7f7fc07fffff803fffff007fffff003fffff001fffff003fffff001fffff801f7f7fc01fffffc01fffffc01fffefe01fffc7e05fff87e03fffc5c07fffc0807f7ff0007ffff0003ffff0005fffe0003ffff00017";
 when "00001010111" => data <= 768x"ffffffffffffc7ffffffc0ff7f7fc07fffff803fffff005fffff003fffff001fffff001fffff001fffff801f7f7fc01fffffc01fffffc01fffefe00fffc7e01fff83e03fffc5c07fffc0807f7ff0007ffff0003ffff0005fffe0003ffff00017";
 when "00001011000" => data <= 768x"ffffefffffffc7ffffffe0ff7f7fc07fffff803fffff001ffffe001fffff001fffff001fffff001fffff800f7f7fc01fffffc00fffffc01fffe7e00fffc7e01fff83e03fffc1c07fffe0803f7f70007ffff0003ffff0001fffe0001ffff0001f";
 when "00001011001" => data <= 768x"ffffe7ffffffc5ffffffe07f7f7fc07fffff803fffff001ffffe001fffff001fffff000fffff001fffff800f7f7fc017ffffc00fffffc01fffe3e00fffc1e017ffc3e03fffc1c05fffe0803f7f70003ffff0003ffff00017ffe0000ffff0001f";
 when "00001011010" => data <= 768x"ffffe3ffffffc17fffffe03f7f7f401fffff003fffff001ffffe001fffff001fffff000fffff000fffff800f7f7f4007ffffc00ffff7c007ffe3e00fffc1e017ffc3e03fffc1c05fffe0803f7f70003ffff0003ffff00017ffe0000ffff0001f";
 when "00001011011" => data <= 768x"ffffe3ffffffc17fffffe03f7f7f401fffff001fffff001ffffe000fffff0017ffff000fffff0007ffff800f7fff4007ffffc00ffff5c007ffe1e00fffc1e017ffe1e01fffc0401ffff0003f7f70001ffff0003ffff00017fff0000ffff00017";
 when "00001011100" => data <= 768x"ffffe1fffffff17fffffe03f7f7f001fffff001fffff001ffffe000fffff0007ffff0007ffff0007ffff80077fff4007ffffc007fff5c007ffe0e007ffc1e017ffe0e01ffff0401ffff8003f7f70001ffff0001ffff0001ffff00003fff01017";
 when "00001011101" => data <= 768x"ffffe1fffffff05fffffc01f7f7f001fffff000fffff0007fffe000fffff0007ffff0007ffff4007ffff80077fffc007ffffc007fff1c007ffe0e007fff17017ffe0e00ffff0401ffff8003f7ff0001ffff8001ffff0001ffff0000bfff01007";
 when "00001011110" => data <= 768x"ffffe0fffffff01fffffc01f7f7f001fffff000fffff0007fffe0007ffff0007ffff0007ffff4007ffff80077f7fc007fffbc003fff0c007ffe0e003fff07017fff0600bfff0401ffff8000f7ff0001ffff8001ffff0001ffff8000bfff01007";
 when "00001011111" => data <= 768x"fffff0fffffff01fffffc00f7f7f001fffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7fc007fffac003fff04007ffe0e003fff07017fff0200bfff44017fff8000f7f740017fff8001ffff0001ffff8000bfff00017";
 when "00001100000" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0017ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7fc007fff8c003fff04007fff06003fff07003fff0200bfffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "00001100001" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0017ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "00001100010" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "00001100011" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007ffff0007ffff0003ffff0007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "00001100100" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007fff70007ffff0003ffff0007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff05011";
 when "00001100101" => data <= 768x"fffff0ffffffd05fffffc00f7f7f001fffff000fffff0007fffe0007fff70007ffff0003ffff0007ffff80037f7f0007fff84003fff04007fff06003fff06003fff82003fffc0007fffc000f7f7c0017fff8001ffff0001ffff8000ffff04011";
 when "00001100110" => data <= 768x"fffff0fffffff05fffff800f7f7f001fffff000fffff0007fffe0007ffff0007ffff0003ffff0007ffff80037f7f0007fff88003fff04007fff06003fff06003fff02003fffc0007fff8000f7ff40017fff8001ffff0001ffff8000ffff04011";
 when "00001100111" => data <= 768x"fffff0fffffff05fffff800f7f7f001fffff000fffff0007fffe0007ffff0007fffe0007ffff0007ffff80037f7f0007fff8c003fff04007ffe06003fff04003fff0200bfff40007fff8000f7f780017fff8001ffff0001ffff8000ff7f04011";
 when "00001101000" => data <= 768x"ffffe0ffffffd05fffff801f7f7f001ffffe000fffff0007fffe000ffffc0007fffe0007ffff0007ffff80037f7f0007fff88003fff04007ffe0e003fff04017fff0600bfff04007fff8000f7f710017fff8001ffff0001ffff8000ffff04011";
 when "00001101001" => data <= 768x"ffffe0ffffffd05fffff801f7f7f001ffffe000ffffc0007fffe000ffffc0007fffe0007ffff0007ffff80077f7f0007fffb8003fff04007ffe0c003fff04017fff0600bfff04017fff8000f7f71001ffff8001ffff0001ffff8000ffff04001";
 when "00001101010" => data <= 768x"ffffc3ffffffc07fffff803f7f7f011ffffe001ffffc001ffffc000ffffc0007fffe0007fffd0007ffff00077f7f0007fffb8007fff1c007ffe0c007fff14017ffe0e00bfff0401ffff8000f7ff1001ffff0001ffff0001ffff0000ffff04011";
 when "00001101011" => data <= 768x"ffff83ffffffc07fffff803f7f7f011ffffe001ffffc001ffffc000ffffc0017fffc000ffffc0007ffff000f7fff0007ffff8007ffd1c007ffe0c007ffc1c017ffe0c00ffff0401ffff8000f7ff0001ffff0001ffff0001ffff0000ffff10011";
 when "00001101100" => data <= 768x"ffff03ffffff807fffff803f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc000fffff000f7f7f0007ffff000fffd5d007ffe1800fffc1d017ffe0c03fffc0401fffe0001f7f70001ffff0003ffff0001ffff0001fff700017";
 when "00001101101" => data <= 768x"ffff02ffffff007fffff803f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc001ffffe000f7fff0017ffff800ffff7901fffe3900fffc11017ff81a03fffc1c01fffc0801f7f70001ffff0003ffff0001fffe0001ffff00017";
 when "00001101110" => data <= 768x"fffe00ffffff007fffff003f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc001ffffe000f7fff001fffff800fffff901fffff980fffd71017ff83a03fffc1c01fff81801f7fc0001fffe0003ffff0001ffff0003ffff00017";
 when "00001101111" => data <= 768x"fff800fffffc007ffffe007f7f7c003ffffc003ffffc001ffff8001ffff8001ffff8000ffffc001ffffe000f7f7f001fffff800fffff101fffff880ffff71017ffaf803fff07c01fff07803f7f07c01fff80803fffc0001fffe0003fff700017";
 when "00001110000" => data <= 768x"ffe001fffff001fffff000ff7ffd007ffff8003ffff0001ffff8003ffff0001ffff0001ffff0001ffff8000f7f7f001fffff001fffff005fffff800fffff1037ffffa03fffffc01fffff800f7f1fc11ffe1f800ffc1fc01ffc0a800ff400001f";
 when "00001110001" => data <= 768x"ffe303ffffc001ffffc000ff7f70017ffff0007ffff0007ffff0003ffff0001ffff0003ffff0001ffff0001f7f75001fffff001fffff101ffffe000ffff7501fffff201fffff401fffff800f7f7f4017ffffc007ffffc017ffbfc003fc17c013";
 when "00001110010" => data <= 768x"ffffe7ffffd541ffffc001ff7fc0017fffe0007ffff0007ffff8003ffff0013ffff0003ffff0001ffff0001f7f70001ffffa001fffff001ffffe000fffff501ffffe581ffffc501ffffee00f7f7f4007ffffe007ffff4007ffffe003ffffc001";
 when "00001110011" => data <= 768x"fffffffffffffdfffffee0ff7f70007ffff0003ffff0005ffffc003ffffc001ffff8001ffffc001ffff8000f7f7c001ffff8000ffffd000fffff000fffff4017fffe080fffff5c07fffe78077f7f5007fffef803fffff001fffff001fffff001";
 when "00001110100" => data <= 768x"ffffffffffffffffffffffff7f7fc51fffff800fffffc007ffff800fffff0007ffff0007ffff0007fffe00037f7f0007ffff0003ffff4007ffffc003fff7c007ffffc003ffffc407ffff8e037f7f1f01ffffbe00ffff7c00fffffc00fffffc00";
 when "00001110101" => data <= 768x"fffffffffffffffffffffe3f7f7f7f17fffffe03fffff401fffff000fffff001ffffe000ffffc000ffffc0007f7fc000fffff000fffff000fffff000fffff000fffff800fffff100fffffb007f7f7701fffff700ffffff00ffffff00fffff700";
 when "00001110110" => data <= 768x"fffffff0fffffff0ffffff807f7f7f00fffffe00fffffc00fffffc00fffffc00fffffc00fffffc00fffffe007f7f7700fffffe00ffffff00fffffe00ffffff40ffffff80ffffffc0ffffff807f7f7fc0ffffff80ffffffc0ffffff80fffff790";
 when "00001110111" => data <= 768x"fffffffffffffff4ffffffe07f7f7f41ffffff80ffffffc0ffffff80ffffffc0ffffffc0ffffffc0ffffffc07f7f7f40ffffffe0ffffffd0ffffffc0ffffff40ffffffc0ffffffc0ffffffc07f7f7f00ffffff00fffffd00fffffe00fffff400";
 when "00001111000" => data <= 768x"fffffffffffffffdfffffff87f7f7f71fffffff0fffffff0fffffff0f7f7fff0fffffff0fffffff0fffffff0757f7f74fa3ffff8f4557c40f0202800f0400000f0200000f5400100ffe002007f500700ffe00200ffc00100ffe00000ffd00100";
 when "00001111001" => data <= 768x"ffff0fffffff57ffffff8fff777f477ffeba03fff50007fffe0003fefd0001f5ff0003f8ff0001f4ff8000f87f400170ff800020ffc00000ffe00000f7701510fff03f80fff47dc0ffffff807f777f00ffffff00ffffff00ffffff00f7f7f700";
 when "00001111010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f5fffffffbffffffd5ffffffbaffffff557fffff23fffffd55fffffe03f7f7f517fffff803fffff407fffff803fffff0037";
 when "00001111011" => data <= 768x"fffbffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00001111100" => data <= 768x"fff03ffffff07ffffff8ffff7f7d7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00001111101" => data <= 768x"fffffffffff07ffffff03fff7ff11f7ffff03ffffff01ffffffc7fffffff7fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00001111110" => data <= 768x"ffffffffffffffffffffffff7f7d7f7ffff81ffffff01ffffff80ffffff01ffffff81ffffffc7fffffffffff7f7fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00001111111" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffff5ffffffc1ffffff41ffffff80ffffff00ffffff80fff7f7c1f7ffffe3fffffff7fffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010000000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff7ffffffe3ffffffc1ffffffc0fff7f7c077ffff807fffffc07fffffc0fffffff5fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010000001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffffffffffffe0fff7f7c077ffff807fffffc07fffff807fffff407fffffe0fffffff5fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010000010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f5f7ffffe0ffffffc07fffffc07fffffc07fffff803fffffc07fffffe0fff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010000011" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7fffffbfffffff1ffffffc07fffffc07fffff803fffffc07fffffc07ff7f7c07ffffff3ffffffffffffffffffffffff7ff";
 when "00010000100" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7fffffffffffff17fffffc07fffffc07fffff803fffffc05fffffc07ff7f7c077fffff0fffffffdfffffffffffffffffff";
 when "00010000101" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffff3ffffffc07fffffc07fffffc07fffff803fffffc07fffffc07ff7f7f177fffff3ffffffffffffffffffffffff7ff";
 when "00010000110" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f177ffffe07fffffc07fffff803fffffc07fffff803fffffc07fffffe0fff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010000111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffff1ffffffe0fff7f74077ffff803fffffc07fffff803fffffc07fffffe0fffffff5fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff7ffffffe0ffffffc07fffff807ff7f70077ffff803fffff407fffffc0ffffff51fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffe3ffffffc17fffff807fffff007fffff807ff7f7107fffff807fffffc07fffffe9fffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001010" => data <= 768x"ffffffffffffffffffffffff7f7fff7ffffffffffffd5ffffffc0ffffff017fffff007fffff007fffff807ff7f70077ffff80ffffffc5ffffffeefffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001011" => data <= 768x"ffffffffffffffffffffffff7f7fff7fffffffffffff5ffffffc0ffffff007fffff807fffff007fffff003ff7f70077ffff80ffffffc1fffffffbffffff7ffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffff7ffffffe1ffffffc07fffff807fffff007fffff803ff7f7003fffff807fffffc07fffffe3fffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001101" => data <= 768x"ffffffffffffffffffffffff7f7fff7fffffffffffffdfffffffbffffffc17fffff803fffff801fffff803ff7f7803fffff803fffffc07fffffe0fffffff5fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001110" => data <= 768x"ffffffffffffffffffffffff7f7fff7ffffffffffffffffffffffffffffd07fffffe03fffffc01fffff803ff7f71017ffff803fffffc01fffffe07ffffff17ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010001111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff57fffffe03fffffc01fffffc01ff7f7c01fffff801fffffc01fffffc03fffff407ffffff2fffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffff83fffffd05fffffc01ff7f7c01fffff801fffffc01fffffc01fffff401ffffff03ffffff57ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffffffffafffffff05fffffe01ff7f7c01fffffc01fffffc01fffffc01fffff401fffffe03ffffff57ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffbfffffff07fffffc03ff7f7c017ffff801fffffc01fffffc01fffff407fffffe03ffffff1dffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffff07fffffc03ff7f7c017ffff803fffffc01fffff803fffffc117ffffe03ffffff47ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010100" => data <= 768x"ffa00000fffd5555ffffffff7f7ffffffffffffffffffffffffffffffff7fff7fffffffffffc07fffffc03ff7f7c037ffff803fffffc01fffff803fffffc07f7fffc07fffffd1fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00010010101" => data <= 768x"20000000d5540000fffc00007f7c0001fffe0000ffff5400fffffe00f7ffff11fffffe03ffff0505fffc06037f740701fff80380fff40741fff80380f7fc0751fffc07f2fffd1fd5fffffffa7f7f7f77ffffffffffffffffffffffffffffffff";
 when "00010010110" => data <= 768x"022bffff0005ffff0007ffff0007ff7f0003ffff0001c17f0000e07f0001c0770001e03e0001f01c0003f80800077800000ff8000007fc000007fc000007fc000003f8000001f000000020000000000000000000000000000000000000000000";
 when "00010010111" => data <= 768x"022bffff0005ffff0007ffff0007ff7f0003ffff0001c17f0000e07f0001c0770001e03e0001f01c0003f80800077800000ff8000007fc000007fc000007fc000003f8000001f000000020000000000000000000000000000000000000000000";
 when "00010011000" => data <= 768x"022bffff0005ffff0007ffff0007ff7f0003ffff0001c17f0000e07f0001c0770001e03e0001f01c0003f80800077800000ff8000007fc000007fc000007fc000003f8000001f000000020000000000000000000000000000000000000000000";
 when "00010011001" => data <= 768x"022bffff0005ffff0007ffff0007ff7f0003ffff0001c17f0000e07f0001c0770001e03e0001f01c0003f80800077800000ff8000007fc000007fc000007fc000003f8000001f000000020000000000000000000000000000000000000000000";
 when "00010011010" => data <= 768x"fffffff007fffff007fffff003f7f7f001fffff0017ffff000ffffc0017f7f4003ffff0007fffc0007fff80017f7100007ff000007ff000003ff800001ff000000f800000050000000000000000000000000000000000000000000000000000";
 when "00010011011" => data <= 768x"3fffffff7fffffffffffffffff7f7f7fffffffffffffffffbfffffff3fffffff3fffffff7fffffdffe8eff0f75007701fa007200fc005000fc000000f4001000f8000000f0000000800000000000000000000000000000000000000000000000";
 when "00010011100" => data <= 768x"f8f80000fdfc0000fffc00007ffc0001fffe0000fffc0005fffe003fffff55ffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff57fff22f00bff00700055003800000111000000000000000000000000000000000000";
 when "00010011101" => data <= 768x"000000000000000000000000140000003e0000001c0000003e0000007f000000ff000000ff400000ffc00a807f417ff4ffeffffcfffffffdffffffffffffffffffffffffffffffffffffffff7f77ffffffe0bffe5fc0057c0600003c00100014";
 when "00010011110" => data <= 768x"80000000c000000080000000500000003000000070000000f8000000f0000000f8000000dd000000e3000000f5715540ffffffe0ffdffff0fffffff8f7fffff5fffffffefffffffdfffffffe7f7fff7dff0ffffeff055fd43a000be010000150";
 when "00010011111" => data <= 768x"e0000000f4000000fe00000075000000ff000000df000000ef800000d7400000ff800000ffc00000ffe800007f770000fff38220ffd55ffdfffffffffffffff7ffffffffffffffffffffffffff7f7f7ffffffffffffdfffffff83fff57f0157f";
 when "00010100000" => data <= 768x"fffe0000ffff4000ffff80007f7f4000ffffa000fff54000ffff8000fff70000ffef8000ffdf8000ffff80007f7f0000ffffe200f7ffff40e7ff8f82d7ff55f79fffffffdfffffffffffffffff7f7f7ffffffffffffffffffffffffffffff7ff";
 when "00010100001" => data <= 768x"03fffff801fffffd00fffff8007f7f50003fff80407ffd40f03ffc00f07fff00f87fe300fc7fc740fe7feff01f7f77700ffffff005fffff003fffff001f7ffff01c3ffef01c7ffd5038fffff071f7f7fbfffffffffffffffffffffff157fffff";
 when "00010100010" => data <= 768x"000fffff0007ffff0007ffff00037f7f0000ffff00007ffd00607ffe0170777101f8fff801f17ff400f8ff88005d7fdd000fffff0007ffdf0003ffff0001f7ff0003efff0005c7ff00070fff00071f7f000e3fff001c7fffea3effffffffffff";
 when "00010100011" => data <= 768x"000fffff0007ffff0003ffff00017f7f00007fff00005fff00000fff001417f7001e0fff001f1ffd001e1ffe001f1f7d0003bffb0001dffd0000ffff00007fff00003fff00005dff000070ff0000717f0000e1ff0001c5ff000187ff000117ff";
 when "00010100100" => data <= 768x"000fffff0007ffff0003ffff00017f7f00003fff00001fff00000fff000117ff000303ff0007c5ff000f83ff0007477f00078ffe0005c7ff00007ffe000077ff00003fff00001fff00000fff00001d7f00001c3f00001c7f0000387f0000717f";
 when "00010100101" => data <= 768x"000fffff0007ffff0003ffff00017f7f00007fff00001fff00001fff000017f7000003ff0001c1ff0007c1ff0007c17f0007c3ff0007c7ff0000e7ff000077ff00003fff00001fff00001fff00001f7f00000fff00000d7f00000c3f00001c1f";
 when "00010100110" => data <= 768x"007ffffe001fffff001fffff00177f7f0003ffff0001ffff00007fff00001fff00001fff000145ff0003c3ff0007c1ff000fc3ff0007c1ff0003e3ff000177ff00003fff00007fff00003fff00001f7f00001fff00001fff00000fff00001c7f";
 when "00010100111" => data <= 768x"007ffffe007fffff003fffff011f7f7f0007ffff0001ffff0000ffff00007ff700003fff00011fff00038fff0007d7ff000fc3ff0007c1ff0007c3ff0001c3f7000067ff000077ff00003fff00007f7f00003fff00001fff00003fff000017ff";
 when "00010101000" => data <= 768x"007fffff005fffff001ffffe00177f7f0003ffff0001ffff0000ffff00007fff00003fff00003fff0001bfff0007df7f0007e3ff0007c1ff0007c3ff0007c3ff0000e3ff000077ff00003fff00007f7f00003fff00001fff00003fff00001f7f";
 when "00010101001" => data <= 768x"003fbfff005fffff001fffff001f7f7f0007ffff0005ffff0001ffff000077ff00007fff00007fff00003fff00015f7f0003ffff0007f7ff0007e3ff0001f3f70001f3ff000077ff00003fff00003f7f00003fff00001fff00003fff00001fff";
 when "00010101010" => data <= 768x"007f07ff007fffff001fffff001f7f7f000ffffe0007ffff0003ffff0001f7ff0000ffff00007fff00003fff00007f7f0001ffff0001ffff0003f7ff0003f7f70001f3ff000177ff00003fff00001f7f00001fff00001fff00001fff00001fff";
 when "00010101011" => data <= 768x"00fe0fff01fd1fff00ffffff007fff7f003ffffe001ffffc000ffffe0007f7ff0003ffff0001ffff00007fff00007f7f0000ffff0001ffff0003ffff0001f7ff0001f3ff0001f7ff00003fff00011f7f00001fff00001fff00000fff00001fff";
 when "00010101100" => data <= 768x"00fe1ff8007c1ffc00783fff017d7f7703fffff301fffff100fffff80077f7ff000fffff0005ffff0001ffff00017f7f00007fff0001ffff0001ffff0001f7ff0003f7ff0001f7ff00003fff00001f7f00000fff00001fff00000fff00001fff";
 when "00010101101" => data <= 768x"00601ff001c05ff401f87ffc01f07f7700f2ffe3015fffc103ffffe003fff7f501ffffff005fffff0007ffff00017f7f0000ffff0001ffff0001ffff0001f7f70003f7ff0001ffff00003ffe00001f7d00001ffc00001ffc00001ffe00001fff";
 when "00010101110" => data <= 768x"0000020000001fc000003ff000007ff400e0ffbf01f5ffc501ffff8001fff7d000fffffe005fffff000fffff00017f770000ffff0001ffff0003efff0003d7f70003ffff00017fff00003fff00001f7500003ffb00001ffd00003fff000017f7";
 when "00010101111" => data <= 768x"000000000000150000003f8000147fc0003efff0001dff5c00ffff000077f700003ffff80017fffd0003ffff00017f770000ffff0001dfff0003cfff0001dfff0001ffff00007fd500003fe600007ff700003fff000077ff000033ff000073ff";
 when "00010110000" => data <= 768x"00000000000000000000000000147f00003c7f80007dff50003ffe00007fff00000fffe00005fff40000fff800017ff00003bffe0007dffd0003bfff00017f1500007f8000007fdd00007fff0000777f000027ff000047ff0000e7ff0001c7f7";
 when "00010110001" => data <= 768x"0000000000000000000000000000140000087e00001d7f00001ffc800017fc000003ff000001ffc00000ffe000017ff00003bff80001dfd40000ff800000775000007ff800005ff000006ff80000477700008ff340011ffdfe83ffff7ff7f7f7";
 when "00010110010" => data <= 768x"000000000000000000000000000000000002380000057c00000ffa000007f0000003ff000001ff000001ff8000017fc00001ffa000007d400000ffc000007fc000005fe00000dff40000bfff75517f77ffffffff5755ffff0380ffff014077f7";
 when "00010110011" => data <= 768x"000000000000000000000000000000000000200000047c00000ff0000007f0000001fe0000017f0000037f00000177000000fb0000007f000000ff80000057500000bfeb7d557fff0fffffff0151ff7f0020ffff000005550000030000000100";
 when "00010110100" => data <= 768x"0000000000000000000000000000000000000000000770000007e8000001f0000000fc0000017c000001fe00000175000000fe0000005f000000bfc015117f770fffffff0555ffff0000ffff0000051700000200000000000000000000000000";
 when "00010110101" => data <= 768x"0000000000000000000000000000000000020000000570000003e8000001f1000000f80000017c000000e000000174000000be0000013d5406817ffe05777ff70020ffff00005c5f000008060000000000000000000000000000000000000000";
 when "00010110110" => data <= 768x"0000000000000000000000000000000000020000000750000003e000000170000000f800000174000000e8000000740000003f0005417f5c02fffffc001175fc000018b800001414000000000000000000000000000000000000000000000000";
 when "00010110111" => data <= 768x"0000000000000000000000000000000000000000000140000003e0000001f0000001f800000150000000f8000001750000007fe00155fff00008fff8000011700000000000000000000000000000000000000000000000000000000000000000";
 when "00010111000" => data <= 768x"0000000000000000000000000000000000000000000140000003e0000001f0000000f0000001d0000000f0000001754000fbffe00015dff0000030e0000010000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111001" => data <= 768x"0000000000000000000000000000000000000000000140000003c000000170000000f0000000d0000000f80000557f40002bffe0000055c000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111010" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000170000000f0000000d0000000f80000557f400000bf800000010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111011" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000170000000e000000050000000fa0000157f00000023800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111100" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000170000000e000000050000000fe0000157f00000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111101" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000170000000e000000050000000fe0000157f00000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111110" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000150000000e000000070000020fe0000157f00000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010111111" => data <= 768x"0000000000000000000000000000000000000000000140000000c000000140000000e000000070000028ff0000157f00000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000000" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000150000000e000000070000028ff0000157700000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000001" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000170000000e000000154000039ff0000157700000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000010" => data <= 768x"00000000000000000000000000000000000000000001c0000003c000000150000000e00000015400003bff0000155700000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000011" => data <= 768x"00000000000000000000000000000000000000000005c0000003c0000001c0000000e00000415400003bff0000015700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000100" => data <= 768x"00000000000000000000000000000000000000000005c0000003c0000001c0000000e00000415400003bff0000015700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000101" => data <= 768x"00000000000000000000000000000000000000000005c0000003c0000001c0000001e00000415400003bff0000015700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000110" => data <= 768x"00000000000000000000000000000000000000000005c0000003c0000001c0000001e00000415400003bff0000115700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011000111" => data <= 768x"0000000000000000000000000000000000000000000540000003c0000001c0000001a00000015400002bfe0000115700000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001000" => data <= 768x"000000000000000000000000000000000000000000054000000380000001c000000180000001d0000028fe0000155f00000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001001" => data <= 768x"000000000000000000000000000000000000000000054000000380000001c0000001e0000001d0000000fe0000157f00000003000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001010" => data <= 768x"000000000000000000000000000000000000000000010000000380000001c0000001e0000001c0000000ea000055ff0000006f000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001011" => data <= 768x"00000000000000000000000000000000000000000000000000038000000140000001e0000001c0000000e0000055ff000000ff000000440000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001100" => data <= 768x"00000000000000000000000000000000000000000000000000038000000140000001e0000001c0000000e000005577000001ff000000450000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001101" => data <= 768x"00000000000000000000000000000000000000000000000000028000000140000001e0000001c0000000e00000557700000bff000000450000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001110" => data <= 768x"00000000000000000000000000000000000000000000000000028000000140000001e0000001c0000000e00000557700000bff000000450000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011001111" => data <= 768x"00000000000000000000000000000000000000000000000000038000000140000001e0000001c0000000e000005577000001ff000000450000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010000" => data <= 768x"000000000000000000000000000000000000000000000000000380000001c0000001e0000001c0000000e00000557f000000ef000000450000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010001" => data <= 768x"00000000000000000000000000000000000000000001400000038000000140000000e0000001c0000000fa0000157f0000002f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010010" => data <= 768x"0000000000000000000000000001000000000000000140000001c000000140000000e000000140000000fa0000157f00000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010011" => data <= 768x"0000000000000000000000000000000000000000000140000001c000000150000000e000000070000008fe0000157700000023000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010100" => data <= 768x"0000000000000000000000000000000000000000000140000000c000000170000000e000000074000038ff0000157700000022000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010101" => data <= 768x"0000000000000000000000000000000000000000000140000000e000000170000000e00000007500000aff8000057700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010110" => data <= 768x"0000000000000000000000000000000000000000000140000000e000000170000000e00000007500000eff8000007700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011010111" => data <= 768x"00000000000000000000000000000000000020000000700000007000000070000000380000005540000effc000015540000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011011000" => data <= 768x"00000000000000000000000000000000000018000000740000003c000000140000001e0000001d50000ebff80001157c000000300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011011001" => data <= 768x"0000000000000000000000000000000000000e0000001d0000000f800000150000000f000000075400028ffe0001577f0000033e0000010400000000000000010000000000000000000000000000000000000000000000000000000000000000";
 when "00011011010" => data <= 768x"000000000000000000000000000001000000060000001f4000000f800000070000000780000007d4000007ff000157ff000023bf0000010500000000000000100000000000000000000000000000000000000000000000000000000000000000";
 when "00011011011" => data <= 768x"00000000000000000000000000000100000003000000170000000fc00000074000000380000005c0000003ff000157ff00003fff000005d500000080000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011011100" => data <= 768x"00000000000000000000000000000000000003000000070000000f80000007c00000038000000740000003e20000077f00003fff000055df00000083000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00011011101" => data <= 768x"00000000000000000000000000000000000000000000070000000e00000017000000078000000740000003800000077c000027fe000057ff000002be000001104000000040000000c000000040000000e0000000c0000000c0000000c0000000";
 when "00011011110" => data <= 768x"00000000000000000000000000000000000000000000040000000e00000017000000070000000500000007000000077100000ff000001ff0000007f00000011000000000c1000000c30000007f000000ff000000ff000000ff000000ff000000";
 when "00011011111" => data <= 768x"00000000000000000000000000000000000000000000040000000c000000150000000e000000040000000e000000074000000fe000001fc000000bc010000100300000007c1000007c1800007f500000fff00000fff00000fff80000fff00000";
 when "00011100000" => data <= 768x"00000000000000000000000000000000000000000000040000000c0000001d0000000e000000040000000e000000074000000fc000001fc000000bc010000100300000007c1000007c1800007f500000fff80000fff00000fff80000fff00000";
 when "00011100001" => data <= 768x"00000000000000000000000000000000000000000000040000000c0000001d0000000e0000000c0000000e000000074000000fc000001fc000000b8010000000300000007c1000007c0800007f500000fff80000fff00000fff80000fff00000";
 when "00011100010" => data <= 768x"00000000000000000000000000000000000000000000040000000c0000001d0000000e0000000c0000000e000000074000001fc000001fc00000028010000000380000007c1000007e0800007f700000fff80000fff00000fff80000fff00000";
 when "00011100011" => data <= 768x"00000000000000000000000000000000000000000000040000000c0000001d0000000e0000000c0000000e80000017c000001fc0000017c00000020010000000380000007c1000007e0800007f700000fff80000fff00000fff80000fff00000";
 when "00011100100" => data <= 768x"00000000000000000000000000000000000000000000040000000c0000001d0000000e0000001d0000000f80000017c000001fc0000017400000000010000000380000007c1c00007e0800007f700000fff80000fffc0000fff80000fff00000";
 when "00011100101" => data <= 768x"00000000000000000000000000000000000000000000040000000c000000150000000e0000001d0000000f8000001fc000003f80000015400000000010000000380000007c1c00003e0800007f700000fff80000fffc0000fff80000fff00000";
 when "00011100110" => data <= 768x"00000000000000000000000000000000000000000000040000001c0000001c0000000c0000001d0000000f8000001fc000003f80000015400000000010000000380000007c0c00003e0800007ff40000fff80000fffc0000fff80000fffc0000";
 when "00011100111" => data <= 768x"000000000000000000000000000000000000000000000c0000001c0000001c0000000c0000001d0000000f8000001fc000001f80000005400000000010000000380000007c0400003e0800007ff40000fff80000fffc0000fff80000fffc0000";
 when "00011101000" => data <= 768x"000000000000000000000000000000000000000000000c0000001c0000001c000000080000001d0000000f8000001fc000001f80000005000000000010000000380000007c0400003e0800007ff40000fff80000fffc0000fff80000fffc0000";
 when "00011101001" => data <= 768x"00000000000000000000000000000000000000000000040000001c0000001c0000000c0000001d0000000f8000001fc000003f80000005000000000010000000380000007c0400003e0c00007ff40000fff80000fffc0000fff80000fffc0000";
 when "00011101010" => data <= 768x"0000000000000000000000000000000000000000000014000000180000001c0000000c0000001d0000000f8000001fc000003f80000015000000000010000000380000007c0400003e0c00007ff40000fff80000fffc0000fffc0000fffc0000";
 when "00011101011" => data <= 768x"0000000000000000000000000000000000000000000004000000180000001c0000001c0000001c0000000f8000001f0000003f80000015000000000010000000380000007c0400003e0c00007ff40000fffc0000fffc0000fffc0000fffc0000";
 when "00011101100" => data <= 768x"0000000000000000000000000000000000000000000000000000080000001c0000001c0000001c0000000e0000001f0000003f80000017400000000010000000380000007c0400003a0400007ff40000fffc0000fffc0000fffc0000fffc0000";
 when "00011101101" => data <= 768x"0000000000000000000000000000000000000000000000000000080000001c0000001c0000001c0000000e0000001f0000003f80000017000000020010000000380000007d0400003a0400007ff40000fffc0000fffc0000fffc0000fffc0000";
 when "00011101110" => data <= 768x"0000000000000000000000000000000000000000000000000000080000001c0000001c0000001c0000000e0000001f0000003f8000001f001000020010000000380000007d0400003b8400007ff40000fffe0000fffc0000fffc0000fffc0000";
 when "00011101111" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001c0000001c0000000e0000001f0000003f8000001f0010000b0010000100380000007d0400003b8600007ff40000fffe0000fffc0000fffe0000fffc0000";
 when "00011110000" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001c0000001c0000001c0000001f0000003f8010001f0010000f8010000100380200007d0400003b8600007ff40000fffe0000fffc0000fffe0000fff40000";
 when "00011110001" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001c0000001c0000001c0000001f0000001f8010001f0010000f8010000100380200007d0400003b8600007ff40000fffe0000fffc0000fffe0000fffc0000";
 when "00011110010" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001c0000001c0000001c0000001f0000003f8010001f001800070010000000380200007d0600003b8200007ff70000fffe0000fffc0000fffe0000fffe0000";
 when "00011110011" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001c0000001c0000001c0000001f0000003f80100017001800020010000000380200007d0600003f8200007ff70000fffe0000fffe0000fffe0000ffff0000";
 when "00011110100" => data <= 768x"00000000000000000000000000000000000000000000000000001800000014000000180000001c0000001e0000001f0000003f80100017001800020010000000380200007d0700003f8200007f7f0000fffe0000ffff0000fffe0000ffff0000";
 when "00011110101" => data <= 768x"0000000000000000000000000000000000000000000010000000180000001c000000180000001c0000001e0000001f0000003f801000170018000000100000003c0200007d0700003f820000777f0000fffe0000ffff0000fffe0000ffff0000";
 when "00011110110" => data <= 768x"0000000000000000000000000000000000000000000010000000180000001c000000180000001c0000001e0001001f0000003f801000170018000000100000003c0200007d0300003d820000777f0000fffe0000ffff0000fffe0000ffff0000";
 when "00011110111" => data <= 768x"0000000000000000000000000000000000000000000010000000180000001c000000180000001c0000001e0001001f0000003f001000150018000000140000003c0200007d0100003d820000777f0000ffff0000ffff0000ffff0000ffff0000";
 when "00011111000" => data <= 768x"0000000000000000000000000000000000000000000010000000380000001c000000180000001c0000001f0000001f0000003f001000150018000000140000003c0300007d0100003da300007f7f0000ffff0000ffff0000ffff0000ffff0000";
 when "00011111001" => data <= 768x"0000000000000000000000000000000000000000000010000000380000001c000000180000001c0000001f0000001f0000003f001000150018000000140000003c8300007d8100003de300007f7f0000ffff0000ffff0000ffff0000ffff0000";
 when "00011111010" => data <= 768x"000000000000000000000000000000000000000000001c0000003e0000001c000000180000001d0000000f8000001fc000003f80100017401800000010000000380000007d0100003d81800075550000ffff0000ffff0000ffff0000ffff0000";
 when "00011111011" => data <= 768x"000000000000000000000000000001000000080000001c0000001e0000001c0000001e0000001f0000000fc000001f5000003fe000001fc000000b80100001003000000074000000f80100007d010000fb018000ff550000ffff8000ffff0000";
 when "00011111100" => data <= 768x"0000000000000000000000000000040000000e0000001f0000000f800000170000000e0000001740000007f00000077100000ff800001ffc00000ff8000005500000000040000000e000000050000000f0000000f0010000f0038000f1010000";
 when "00011111101" => data <= 768x"000000000000000000000200000007000000070000001fc000000fc00000070000000f0000001754000003fc000007ff000007ff00001fff00000fff00001777000002fa000004400000000000000000800000000000000080000000c0000000";
 when "00011111110" => data <= 768x"00000000000001400000018000000340000007e000001ff0000003f0000007f000000fc000001dd5000003ff000001ff000003ff000005ff00000fff000017ff00000fff0000057f000001bb0000011100000000000000000000000000000000";
 when "00011111111" => data <= 768x"00000060000000f0000000e0000005f500000ffe000005fc000001fe000001f400001bf000001df5000008ff0000117f000000ff0000047f000000ff000001ff000003ff000007ff000007ff000007ff000000e7000000470000004600000040";
 when "00100000000" => data <= 768x"0000003e0000007f000001ff000007ff000003ff0000007f0000007f0000017f000039ff00005fff00002eff0000103f0000003f0000001f0000001f000000170000003f0000007f000000ff0000017f000003ff000001ff000001ff000001ff";
 when "00100000001" => data <= 768x"000000ff000001ff000003ff0000015f0000000f000000070000000f000000770000707f0001ddff0001cfff0001475700004007000040070000000700000007000000030000000100000003000001030000000300000047000000ef00000077";
 when "00100000010" => data <= 768x"000001ff0000007f0000002000000000000000000000000000000000000000170003803f0007d07f000ff8ff001d7fff000a1fff0007055500020000001300000002000000000000000000000000000000000000000000000000000000000000";
 when "00100000011" => data <= 768x"000000ff0000007d0000000000000000000000000000000000000007000000070003801f0007f07f000ffeff00153fff001a1fff0006054500060000000600000002000000000000000000000000000000000000000000000000000000000000";
 when "00100000100" => data <= 768x"0000003f000000550000000000000001000000000000000000000003000000070003e00f0007f45f000ffeff001d1fff001a0fff001707c500060000000700000002000000050000000000000000000000000000000000000000000000000000";
 when "00100000101" => data <= 768x"0000003f000000140000000000000000000000000000000100000003000000030000e0070005f41f0007fe7f00071f7f000f0fff000507f500030280000100000003000000010000000000000000000000000000000000000000000000000000";
 when "00100000110" => data <= 768x"0000000b000000000000000000000000000000000000000000000000000000010000f0030001fc070003ff3f00075f7f00078fff0005c7fd000383e000010000000180000001c000000000000000000000000000000000000000000000000000";
 when "00100000111" => data <= 768x"00000002000000000000000000000000000000000000000000000000000050010000f8030001fd070003ff9f000757ff000787ff0005c5fd0002c0e80001c0000000c0000000c000000080000000000000000000000000000000000000000000";
 when "00100001000" => data <= 768x"00000000000000000000000000000000000000000000000000000000000050010000f8030005ff470007ffff0017477f000f83ff0005c1fd0000c0e80001c0000000c0000000c000000080000000000000000000000000000000000000000000";
 when "00100001001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000017000000ffe03001fdfd7001ecfff0015077f000003ff0001017d0003800000018000000180000001c0000001c0000001000000000000000000000000000000000000";
 when "00100001010" => data <= 768x"000000000000000000000000000000000000000000000000000000000017f500003fffa100145ff700080fff0000057f000000ff0000007f000000000000000000020000000700000003000000030000000380000001c0000000800000000000";
 when "00100001011" => data <= 768x"00000000000000000000000000177551003ffffb001d7fff000ccfff001445ff000000ff000000550000000000000000000000000000000000000000000000000000000000040000000e00000007000000030000000700000002000000000000";
 when "00100001100" => data <= 768x"000c60ff0004405500000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080000001c000000180000001c0000000e00000007000000000000000000000000000000000000";
 when "00100001101" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000300000001c0000001e0000001700000006000000040000000000000000000000000000000000000000000000000000";
 when "00100001110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000006000000070000003e0000007d000000200000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00100001111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000180000001c0000000c0000001c000000180000001c000000000000001000000000000000000000000000000000000000000000000000000000000000000000";
 when "00100010000" => data <= 768x"00000000000000000000000000000000000000000000000000080000001c000000180000000c0000000e000000070000000600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00100010001" => data <= 768x"00000000000000000000000000000000000000000000000000080000001c0000003f8000000700000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00100010010" => data <= 768x"00000000000000000000000000000000000000000001c000000f8000001f0000000c000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000050000000e800000075000000";
 when "00100010011" => data <= 768x"fff80000fff54000fffe80007f7f5000fffe2000fffc7500fffcfe00f7f1f750fffeffe0ffffffd4fffffffe7f7f7f7dfffffffffffffffffffffffff7fff7f7ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100010100" => data <= 768x"fffffffffffd7ffffffc7fff7f7c7f7ffffe3fffffff1fffffff1fffffff7fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100010101" => data <= 768x"fffffffffffd77fffffe07ff7f7c077fffffa7ffffffd7ffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100010110" => data <= 768x"ffffe3ffffffc5ffffff0fff7f7f1f7fffff3fffffffdffffffffffffffff7ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100010111" => data <= 768x"ffffe3ffffffc7ffffffe3ff7f7f437fffffe7fffffff7ffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100011000" => data <= 768x"fffff03ffffffc7ffffffc7f7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100011001" => data <= 768x"ffff83ffffffc7ffffffc7ff7f7fd7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100011010" => data <= 768x"ffffe0fffffff0fffffff8ff7f7f707ffffff83ffffffc5ffffff8fffffff5ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100011011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffdfffffff9f7f7f571fffffa20fffff541fffff800fffff0117ffff80afffff55dfffffafff7f7f5f7fffffffffffffffffffffffffffffffff";
 when "00100011100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7f7ffffffffffffd57fffffc07f7f7fc07fffffe07ffffff07ffffff0fffffff17ffffff0fffffff1ffffffe0ff7f7f417fffffe0ffffffd5fffffffbfffffff7ff";
 when "00100011101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffd7ffffffc3ffffffc1ffffff81ffffff017fffffe07ff7f7f017fffff80ffffffc1ffffffe0fffffff37fffffffffffffffffffffffff7f7f7ffffffffffffffffffffffffffffffff7ff";
 when "00100011110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7f7ffffe033ffffc005ffffe001ff7f4511ffffc783ffffdfd7ffffffffffff77ffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100011111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff77ffffff80fffffd007ffffc007ff7fc1577fff87ffffffc7ffffff8fffffffdfffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100100000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff57fffffe83fffffc07fffffc07fff7fc77f7fff8fffffff1fffffff0ffffff717ffffff1fffffffdfffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100100001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffff7fdffffffe0ffffff01ffffff83ffff7f177f7fff1fffffff1ffffffe1ffffff71ffffffe3ffffffc1ffffffebfffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00100100010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffeffffff7c7ffffffc3ffffffc7fffffe8fffff7d1f7f7fff1fffffff1ffffffe3ffffff717fffffe3ffffffc7ffffffc3fffff7d3f7f7ffd3ffffffd7fffffffffffffffffffff";
 when "00100100011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffff71ffffffe1fffffff1ffffffe1fffff7c1f7f7ff83ffffff45ffffffe3ffffffc37fffffe3ffffffc7ffffffc3fffff7c3f7f7ff83ffffffd7ffffffd7fffffff7fffff";
 when "00100100100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffefffffffc77fffffc7ffffffc7ffffffc3fffff7c3f7f7ff83ffffff07ffffff87ffffff47ffffff87ffffffc7ffffff87fffff787f7f7ff83ffffff17ffffffb7ffffff77fffff";
 when "00100100101" => data <= 768x"ffffffffffffffffffffffffff7f7f7ffffffffffffffffff8fffffff07ffffff8fffffffc7ffffff87fffff717f7f7ff8fffffff07ffffff0fffffff07ffffff87ffffff07ffffff87fffff717f7f7ff83ffffff17ffffffb7fffffff7fffff";
 when "00100100110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffdfffffff8fffffff077fffff8fffffff07ffffff07fffff707f7f7ff0fffffff1ffffffe0fffffff077fffff8fffffff07ffffff87fffff707f7f7ff87ffffff07ffffffa7ffffff177ffff";
 when "00100100111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffff5fffffff0fffffff077fffff8fffffff07ffffff03fffff717f7f7ff0fffffff07fffffe0fffffff07ffffff8fffffff07ffffff87fffff707f7f7ff87ffffff07ffffff03ffffff17fffff";
 when "00100101000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ff8fffffff07ffffff87ffffff077fffff83ffffff07ffffff03fffff707f7f7ff07ffffff07fffffe07ffffff077fffff87ffffff07ffffff87fffff707f7f7ff83ffffff07ffffff83ffffff17fffff";
 when "00100101001" => data <= 768x"ffffffffffffffffffffffff7d7f7f7ff83ffffff01ffffff83fffff7c77fffff83ffffff01ffffff81fffff705f7f7ff03ffffff07fffffe03ffffff47ffffff83ffffffc1ffffff83fffff711f7f7ff83ffffff01ffffff81ffffff11fffff";
 when "00100101010" => data <= 768x"ffffffffffffffffffffffff7d3f7f7ff83ffffffc1ffffffc3fffff7c1ffffffc0ffffffc1ffffff80fffff7c1f7f7ff83ffffff01ffffff01ffffff41ffffffc1ffffffc1ffffffc1fffff7c1f7f7ff81ffffffc1ffffff80ffffff11fffff";
 when "00100101011" => data <= 768x"ffffffffffffffffffbfffff7c1f7f7ffc1ffffffc1ffffffe1ffffff417fffffc0ffffffc0ffffffc0ffffffc177f7ff81ffffff01ffffff80ffffff41ffffffe0ffffffc1ffffffc0fffff7c1f7f7ff80ffffffc0ffffff80ffffffc07ffff";
 when "00100101100" => data <= 768x"ffffffffffffffffffbfffff7d1f7f7ffc1ffffffc1ffffffe0fffffff17fffffe07fffffc07fffffe07ffff7c077f7ffc0ffffffc07fffff80ffffffd07fffffe0ffffffc07fffffe0fffff7c077f7ffc07fffffc07fffffc07fffffc07ffff";
 when "00100101101" => data <= 768x"ffffffffffffffffffffffff7f1f7f7ffe0fffffff07ffffff0fffffff07ffffff03ffffff07fffffe03ffff7f077f7ffe07fffffc07fffffc07fffff507ffffff07ffffff07fffffe07ffffff077f7ffe03fffffc07fffffc03fffffc07ffff";
 when "00100101110" => data <= 768x"ffffffffffffffffffcfffff7f077f7fff07ffffff07ffffff87ffff7f07ffffff81ffffff01ffffff83ffff7f017f7fff03ffffff07fffffe03fffff703ffffff83ffffff05ffffff03ffffff037f7fff03ffffff01fffffe03fffff701ffff";
 when "00100101111" => data <= 768x"ffffffffffffffffffe7ffff7f437f7fff83ffffffc3ffffffc3fffff7c1ffffff80ffffffc1ffffff80ffff7fc1ff7fff83ffffff01ffffff01ffffff41ffffff81ffffffc1ffffff81ffff7f01ff7fff81ffffff01ffffff01ffffff01ffff";
 when "00100110000" => data <= 768x"fffffffffff7ffffffe3ffff7fc1ff7fffc1ffffffc1ffffffe0fffff7f07fffffe03fffffc07fffffe0ffff7f417f7fff80ffffff00ffffff80ffffff51ffffffe0ffffffc0ffffffe0ffffffc07f7fffc0ffffffc07fffffc0ffffffc077ff";
 when "00100110001" => data <= 768x"fffffffffffdfffffff8ffff7f717f7fffe07ffffff07ffffff0fffff7f077fffff03ffffff01fffffe03fff7f707f7fffe07fffffc07fffffc07fffffd07ffffff07ffffff07fffffe07fff7f707f7fffe07fffffe07fffffe07fffffe07fff";
 when "00100110010" => data <= 768x"fffffffffffffffffffeffff7f707f7ffff03ffffff07ffffff87ffff7f41ffffff81ffffff01ffffff81fff7ff11f7ffff03ffffff05ffffff03ffffff07ffffff03ffffff07ffffff03fff7f707f7ffff03ffffff01fffffe03ffffff01fff";
 when "00100110011" => data <= 768x"fffffffffffffffffffe7fff7f707f7ffff83ffffffc5ffffffc3ffff7fc1ffffff80ffffffc1ffffff80fff7f7c1f7ffff83ffffffc7ffffff83ffffff07ffffff83ffffff01ffffff83ffffff01f7ffff03ffffff01ffffff01ffffff01fff";
 when "00100110100" => data <= 768x"fffffffffffffffffffebfff7f7c1f7ffff81ffffffc1ffffffc3ffff7fc17fffffc07fffffc07fffffc0fff7f7c177ffff81ffffffc1ffffff83ffffffc17fffff83ffffffc1ffffff81ffffff01f7ffff81ffffff01ffffff80ffffff017ff";
 when "00100110101" => data <= 768x"ffffffffffffffffffffbfff7f7d1f7ffffe0ffffffc0ffffffe1ffff7f617fffffe07fffffc07fffffe07ff7f7c077ffffc07fffffc07fffffc1ffffffc17fffffc1ffffffc1ffffffc0ffffffc1f7ffff80ffffffc07fffff80ffffffc07ff";
 when "00100110110" => data <= 768x"ffffffffffffffffffffffff7f7f1f7ffffe0fffffff07fffffe0ffff7f717fffffe03ffffff07fffffe07ff7ff7017ffffe03fffffc07fffffe0ffffffc1ffffffe0ffffffc1ffffffc0fff7f7c077ffffe07fffffc07fffffc07fffffc07ff";
 when "00100110111" => data <= 768x"ffffffffffffffffffffffff7f7f077ffffe07ffffff07ffffff0ffff7ff17ffffff03ffffff05fffffe00ff7fff017ffffe0bffffff07fffffe0fffffff17fffffe0ffffffc07fffffe07ff7f7e077ffffe07fffffc07fffffe03fffffc03ff";
 when "00100111000" => data <= 768x"ffffffffffffffffffffafff7f7f077fffff07ffffff07ffffff0ffff7ff07ffffff03ffffff01fffffe03ff7f7f037ffffe07ffffff07fffffe0fffffff07fffffe0fffffff07fffffe07ff7f7f077ffffe03fffffe07fffffe03ffffff03ff";
 when "00100111001" => data <= 768x"ffffffffffffffffffff8fff7f7f077ffffe07ffffff07ffffff0ffff7ff07fffffe03fffffc01fffffe03ff7f77037ffffe0fffffff07fffffe0fffffff07fffffe07ffffff07fffffe07ff7f7f077ffffe03ffffff07fffffe03ffffff07ff";
 when "00100111010" => data <= 768x"ffffffffffffffffffffafff7f7f177ffffe07fffffc07fffffe0ffff7f507fffff003fffff001fffff803ff7f7f037ffffe03fffffc07fffffe07fffffe07fffffe07ffffff07fffffe07ff7f7f077ffffe03ffffff07fffffe03ffffff03ff";
 when "00100111011" => data <= 768x"ffffffffffffffffffff8fff7f7f077ffffe03fffffc07fffffe0ffff7f707ffffe203ffffc001ffffe003ff7f77017ffffe03fffffc07fffffe07ffffff07fffffe03ffffff07fffffe03ff7f7f077fffff03ffffff01fffffe03ffffff01ff";
 when "00100111100" => data <= 768x"ffffffffffffffffffff8fff7f7f077ffffe03ffffff07ffffff07fff7f707f7ffe201ffffc001ffff8001ff7fd701ffffff01ffffff05ffffff03ffffff03ffffff83ffffff01ffffff03ff7f7f017fffff03ffffff01fffffe01fffff701ff";
 when "00100111101" => data <= 768x"ffffffffffffdfffffff8fff7f7f077ffffe03ffffff07ffffff07fff7ff07f7ffce01ffffc401ffff8000ff7f1501ffffbf01ffffff05ffffff83ffffff03ffffff83ffffff01ffffff83ff7f7f01ffffff01ffffff01fffffe01fffff701ff";
 when "00100111110" => data <= 768x"ffffffffffffffffffffe7ff7f7f077ffffe03ffffff01ffffff03fff7ff07f7ffbf03ffffc400ffff8000ff7f0101ffffbf01ffffff41fffffe03ffffff037fffff83ffffff81ffffff81ff7f7f01ffffff01ffffff01ffffff01ffffff01ff";
 when "00100111111" => data <= 768x"fffffffffffff7ffffffc7ff7f7f077ffffe03ffffff01ffffff03fff7ff03f7ffff81ffff14007fff0000ff7f0101ffff3e00ffffff01fffffe83fffff711ffffff83ffffff01ffffff81ff7f7f01ffffff01ffffff01ffffff01fffff701ff";
 when "00101000000" => data <= 768x"ffffffffffffd7ffffff87ff7f7f017ffffe03fffffe07ffffff03fff7ff03ffffff03fffd5401fffc0000ff7c0101fffe2e01fffdfd01fffffe01fffffd01ffffff03ffffff01ffffff03ff7f7f01ffffff03ffffff01fffffe01fffff401ff";
 when "00101000001" => data <= 768x"ffffffffffffc7ffffff03ff7f7f037ffffe03fffffc07fffffe03ffff7f03ffffff03fffd7c01fffc0000ff7e00017ffe2e01ffff7c01fffffe00fffff701fffffe01fffffe01fffffe01ff7f7f017ffffe03fffffc01fffffe03fffffc01ff";
 when "00101000010" => data <= 768x"ffffffffffffdfffffff87ffff7f077ffffe03fffffc01fffffe03ffffff0177ffff03fffffd41ffffa800ff7f00017fff8201ffffde01fffffe00ffffff017ffffe00ffffff01fffffe00ff7f7f017ffffe00ffffff01fffffe03ffffff03ff";
 when "00101000011" => data <= 768x"ffffffffffffdfffffffefffffff477fffff03ffffff01fffffe01ffffff01f7ffff81ffffff41ffffff80ff7f75007fffe000fffff101fffffe00ffff7f007fffff007fffff007fffff007f7f7f007fffff007fffff007ffffe02ffffff03ff";
 when "00101000100" => data <= 768x"ffffffffffffdfffffffcfffffff017fffff01ffffff01fffffe01ffffff017fffff80ffffff81ffffff80ff7f7f007fffff00fffffc007ffff8007ffff1007fffff003fffff007ffffe003f7f7f007fffff003fffff005ffffe003fffff0377";
 when "00101000101" => data <= 768x"ffffffffffffdfffffff83ffffff017fffff00ffffff01fffffe00fffff7007fffff80ffffffc0ffffff80ff7f7f007fffff80ffffff007fffff007fffff007ffffe003ffffc007ffffe003f7f7f003ffffe003fffff005fffff003fffff007f";
 when "00101000110" => data <= 768x"ffffffffffffdfffffffcbff7f7f017fffff80ffffff007ffffe00fffff7007fffff807fffffc07fffff80ff7f7fc07fffff807fffffc07fffff807fffff007fffff003fffff007fffff003f7f7f003fffff003fffff007fffff007fffff007f";
 when "00101000111" => data <= 768x"ffffffffffffffffffffffff7f7fc57fffff80ffffff007fffff80fffff70077ffff807fffffc07fffffc07f7f7fc07fffffc07fffffc07fffff807fffff0077ffff007fffff007fffff803f7f7f007fffff003fffff007ffffe007fffff0077";
 when "00101001000" => data <= 768x"ffffffffffffffffffffffff7f7f41ffffff80ffffff007fffff80fffff70077ffff807fffffc07fffffc0ff7f7fc07fffffc07fffffc07fffff807fffff0077ffff003fffff007ffffe003f7f7f0077fffe003ffffc007ffffe007ffff5007f";
 when "00101001001" => data <= 768x"ffffffffffffffffffffffff7f7f41ffffff01ffffff01ffffff00ffffff0177ffff80ffffffc07fffffc0ff7f7fc07fffff80ffffffc07fffff807ffff7007fffff003fffff007ffffe003f7f7d003ffff8003ffffc007ffff8007ffff7007f";
 when "00101001010" => data <= 768x"ffffffffffffffffffffffff7f7f077fffff01ffffff01ffffff01fffffd01f7ffff00ffffffc0ffffff80ff7f7f417fffff80ffffff807fffff807ffff7107ffffe003ffffc007ffff8003f7f71003ffff0003ffff5007fffec003ffff50077";
 when "00101001011" => data <= 768x"ffffffffffffffffffffffff7f7f577fffff03ffffff01ffffff01fffffd01ffffff00ffffff01ffffff80ff7f7f017fffff80ffffff007ffffe007ffffc007ffff8003ffff0007fffe0803f7fc1003fffe3003fffd7001fffff003fffff003f";
 when "00101001100" => data <= 768x"ffffffffffffffffffffffff7f7f577fffff81ffffff01ffffff00ffffff01ffffff00ffffffc1ffffff80ff7f7fc1ffffff80ffffff00fffff800fffff0007fffc0007fffc1007fff83803f7f67007fffef003fffff007fffff003ff7ff0077";
 when "00101001101" => data <= 768x"ffffffffffffffffffffcfff7f7f41ffffff80ffffff007fffff00fffff70077ffff80ffffffc1ffffffc0ff7f7f41fffffe00ffffd0007fff8000ffff01017fff8300ffff47007fffde007f7fff007fffff00ffffff007fffff80ffffff0077";
 when "00101001110" => data <= 768x"ffffffffffffdfffffffc3ff7f7fc1ffffff80ffffff007ffffe00fffff70077ffff807fffffc0ffffffc0ff7ff5017fff8000ffff00007fff0380fff75700f7ff9f00ffffff007ffffe00ff7f7f017fffff80ffffff01ffffff80ffffff01f7";
 when "00101001111" => data <= 768x"ffffffffffffffffffffefff7f7fc1ffffff80ffffff407fffff007fffff407fffffc07fffffc07fffebc0ff7f00017ffe0000ffffc4007fffcf80ffffdf0077ffff00ffffff007fffff80ff7f7f017fffff80ffffff81ffffff80ffffff01f7";
 when "00101010000" => data <= 768x"ffffffffffffffffffffefff7f7ff17fffffc07fffffc07fffff803fffffc07fffffc03ffd45c07fffe0807f7fc0017fffe0007fffd7407fffff807ffff7007fffff007fffff007fffff807f7f7f007fffff007fffff007fffff80ffffff0177";
 when "00101010001" => data <= 768x"fffffffffffff7fffffff3ff7f7ff17fffffe03fff7f401fffbf803fffc7c037ffe1e03fffe0405fffe0003f7fd5017fffff003fffffc07fffff803fffff007fffff003fffff007fffff803f7f7f003ffffe003ffffd007fffff803fffff017f";
 when "00101010010" => data <= 768x"fffffffffffffdfffffff0ff7fdf707fffdfa03fffc7c01fffe3e01ffff15017ffe0603ffff0401fffec003f7f7f013fffff803fffffc01fffff803fffff001fffff003fffff001fffff001f7f7f001fffff001fffff001fffff001fffff001f";
 when "00101010011" => data <= 768x"fffffffffff7fdffffeff87f7f77701fffe3801ffff5c01ffff8e01ff7f0701ffff0203ffff4001fffff003f7f7f401fffff803fffffc01fffff803fffff001fffff001fffff001fffff000f7f7f001fffff000fffff0007ffff000fffff0007";
 when "00101010100" => data <= 768x"ffffffffffffff7ffffffe7f7f73f41ffff3e01ffff1c00ffff9e00ffffd7007fff8700ffffc501ffff8001f7f77011fffff801fffffc01fffff801ffff7001fffff001fffff001fffff000f7f7f0117ffff000fffff0007ffff800fffff0007";
 when "00101010101" => data <= 768x"ffffffffffffff7ffffffc3f7f7ff01fffffe00fffffc007ffffc00ffffdd007fff8e007fff9f007fff8f0077f7d7007fffc6007fffc4007fff80007fff40007fffe0003ffff0007ffff00037f7f0003fffe0003fffd0001ffff0003ffff0101";
 when "00101010110" => data <= 768x"ffffff3ffffff41ffffff0077f7ff007ffffe003ffff4007ffff8003fff74003ffffe003fffff001fffff0017f7f5001fffe3000fffc7000fffc6000fffc7000fffe0000fffc0000fffe00007f7c0000fffc0000fffd0000ffff8000fff7c000";
 when "00101010111" => data <= 768x"fffffe01fffffc00fffff8007f7f7000ffff8000ffffc000ffff8000ffffc000ffffe000fffff000fffff0007f7f7000ffffb000fffd7400fff86000fff07000fff8f000fff87000fff820007f7c0000fffe0000fffc0000fffe0000fff40000";
 when "00101011000" => data <= 768x"fffffe00fffffc00fffff8007f7f7000fffff000ffffc000ffff8000ffff0000ffff8000ffffc000ffefe0007ff77000fff7f000ffd7f000ffc3f200ffc3f100ffe3f200ffc1f000ffe1e0007f714000fff80000fffc0000fff80000fff40000";
 when "00101011001" => data <= 768x"fffffe03fffffc00fffff0007f7f7100fffff000ffffd000ffffc000ffff0000ffff0000ffdfc000ffefc0007ff77000ffe7f000ffc7f000ff83f000ffc3f000ffe3f000ffc1f000ffe1e0007f714000fff80000fffc0000fff80000fff00000";
 when "00101011010" => data <= 768x"fffff803fffff001ffffe0007f7f7000ffffe000ffffc000ffff8000ffff0000ffff0000ffff4000fffee0007f7df000fff1e000ffc1f000ffe1e000fff1f000ffe3e000fff1f000fff0e0007f704000fff80000fffc0000fff80000fff00000";
 when "00101011011" => data <= 768x"fffff803fffff001ffffe0007f7fc000ffff8000ffff0000fffe0000ffff0000ffff8000fffdc000fffde0007f7dc000ffe3e000ffc1c000ffc3e000ffc1c400ffe3e000ffc1c000ffe1e0007ff14000fff80000fffc0000fff80000fff00000";
 when "00101011100" => data <= 768x"fffff80ffffff005ffffe0017f7fc001ffff8000ffff0000fffe0000ffff0001ffff8000ffdfc000ffcfc0007f5f4000ffefe000ffc7c000ff87c800ff07c401ff83c000ffc5c001ffe1c0007f714001fff00000fffc0001fff80000fff00001";
 when "00101011101" => data <= 768x"ffffff0ffffff405fffff0017f7f7001ffffe000ffffc000ffff8000fff70000ffff0000ffffc000ffbfe0007fdf4000ffcfe000ffc7c000ff87c000ff07c400ff83c400ffc5c000ffe180007f710001fff00000fffc0000fff80000fff00000";
 when "00101011110" => data <= 768x"fffff801fffff001ffffe0007f7f7000ffffe000ffffc000ffff8000fff70000ffff8000fffdc000fff9e0007f7df000ffe3e000ffc1f000ffc3e000ffc3f600ffe3e200ffc1c000ffe0c0007ff10000fff80000fffc0000fffc0000fffc0000";
 when "00101011111" => data <= 768x"fffff800fffff000fffff0007f7f7000ffffe000ffff4000ffff0000ffff0000ffffc000ffff5000fffef0007f75f000ffe1f000ffc1f000ffe1f200fff1f100ffe3f200fff1f000fff8e0007f704000fff80000fffc0000fffe0000fffc0000";
 when "00101100000" => data <= 768x"fffffc00fffffc00fffff8007f7ff000fffff000ffffc000ffff8000ffff0000ffffe000ffdff000ffeff8007f5ffc00ffaff800ff07fc00ff07f880ff077c00ff83f880ffc1fc00ffe1f8007f715000fff00000fffc0000fffc0000fff60000";
 when "00101100001" => data <= 768x"ffffff00ffffff00fffffe007f7f7700fffffe00fffff400ffffe000fffff000ffffe000ff7ffc00ff3ffe007fdf7700ffcfff00ffc7ff00ff87ff00ff07ff10ff83ff10ffc1ff10ffe0ff007f707f00fff03800fffc0000fffc0000fffc0000";
 when "00101100010" => data <= 768x"ffffffe0ffffffc0ffffffe07f7f7fc0ffffff00fffffc00fffffc00fffdfd00fffeff00fffc7fc0fffeffe07f7c7f70fff0fff0ffc07ff0ffc07ff0ffc077f1ffe07ff0fff07ff0fff07ff07f7037f0fff81fe0fffc1f40fffe0000fff70000";
 when "00101100011" => data <= 768x"ffffff80ffffffc0ffffff807f7f7f00ffffff80fffffdc0fffffde0fffff1f0fffffbfafffff7fffffe27ff7f7c07fffff807fffffc07fffff80ffffffc17fffff80ffffffc1ffffff80fff7f7d1f7ffffc07fffffc07fcffff03f8ffff1151";
 when "00101100100" => data <= 768x"fffffff8fffffffcfffffffe7f7fff7fffff3fffffff1fffffff3fffffff1fffffff3fffffff1fffffff3fff7f711f7ffff01fffffc01fffffe00fffffc01fffffe00ffffff01ffffff00fff7f70177ffff807fffffc07fffffc03ffffff01ff";
 when "00101100101" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffff5fffffff9fffffff1fffffffc7ffffffc7ffffffe3ffff7f717f7fffe07fffffc07fffff803fffff101fffff003fffff001fffff001fff7f401f7fffe00ffffff007fffff803fffff001ff";
 when "00101100110" => data <= 768x"ffffffffffffffffffffffff7f757f7ffff8fffffff47ffffff87ffffff47ffffffe3ffffffc7ffffffe3fff7f751f7ffff00fffffc00fffff800fffffc007ffff8007ffffc007ffffe00fff7ff0077ffff00ffffff007fffff803fffffc01ff";
 when "00101100111" => data <= 768x"ffffffffffffffffffffffff7f7f7f5fffffff9fffffff1fffffff1ffffff73ffffffe3ffffff47fffff807f7f7d007ffff8007ffffc007ffffc007ffffc007ffffc00fffffc00fffffc00ff7f7c01fffffe03fffffc01fffffe007ffff7007f";
 when "00101101000" => data <= 768x"ffffffffffffffffffffffff7f7fd77fffff8fffffffd7ffffff8fffffffd7ffffff8ffffffd57fffff80fff7f71077fffe007ffffc007ffffc007ffffc007fffff007fffff007fffff00fff7f70077ffff803fffffc01fffffc00fffff4017f";
 when "00101101001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffcfffffffcffffffff7ffffffe3fffffff1fffffff9ffff7f517f7fff807fffff407fffff003fffff003fffff003fffff001fffff803fff7fc01f7fffe00ffffff007fffff001fffff0007f";
 when "00101101010" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffff3fffffff1ffff7ff8fffffffc7ffffffe3ffff7f71ff7fffe07fffffc07fffff803fffff001fffff801fffff001fffff001fff7f401f7fffe007fffff001fffff800fffffc0077";
 when "00101101011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffff9fffffffd7ffffffe3fffffff1fffffff83fff7f701f7ffff00fffffc007ffffc007ffffc007ffffc007ffffc007ffffe003ff7ff0017ffff8003ffffc001ffffe000ffff70011";
 when "00101101100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffd7fff7ffe3fffffff1fffffff8efff7f7c177ffff813fffff401fffff803fffff001fffff001fffff001fffff800ff7f7c005fffff000fffff0005ffffc000ffffd000";
 when "00101101101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7f7ffffffffffdfffffffcfffff7f47df7ffff38ffffff14ffffff00ffffff007ffffe007ffffc007ffffe003ff7f70017ffff00062fffc0000fffe0000ffff0000";
 when "00101101110" => data <= 768x"ffffffe0ffffffc0ffffff807f7f7f00ffffff80ffffffd0fffffff8fffff7fcfffffff8fffffffcfffffffe7fdf7f7fffcefbfeffc67174ffc27060ffc07000ffc00000ffc00000ffc000007f400000ffe00000fff40000fffe0000fff75000";
 when "00101101111" => data <= 768x"fffffc00fffffc00fffffc007f7f7d00fffff000fffff000ffffe000fff7fc00fffffe00fffffc00fffffe007fff7f41fffe7f00fff45c00ffe01800fff01000ffe00000ffc00000ffe000007ff00000fffe0000ffff4000ffffe000fff7f000";
 when "00101110000" => data <= 768x"fffff000ffffc000ffffe0007f7f4001ffffe001ffffc005ffff8007ffff4007ffffe007ffffc007ffffe00f7f77741ffff3f00fffc1c007ffc08003ff001001ff000001fd5c0000fffc00027f7f0007ffff0007ffff4007ffffe007fffff007";
 when "00101110001" => data <= 768x"fffffbefffffc047ffff80077f7f0107ffff000fffff005ffffe003fffff003fffff803fffff007fffff803f7fdfd17fff8f80ffff05001fff00001ffd00001ff8200000fd740010fffc00387f7c007cfffe003fffffc07fffff807fffff0077";
 when "00101110010" => data <= 768x"ffffffffffffd77fffff023f7f7f001ffffe003ffffc007ffffe00bff7fc017ffffe00ffffff01fffffe00ff7f7f477fff3f03fffc1c01fffc0c00fff0000054e0800000fdd001c0fff800e07f790177fff801ffffff05fffffe03fffffc01ff";
 when "00101110011" => data <= 768x"fffffffffffffffffffe0eff7f7c017ffffc007ffffc017ffffc00fffff001fffff803fffffc07fffffc03ff7fff177ffcfe03fffc7c01fdf81803f8f0000150c3000200d7740700fff803db7f70077ffffc07fffffc07fffff80ffffffc07ff";
 when "00101110100" => data <= 768x"fffffffffffffffffffc3bff7f78117ffff801fffff001fffff803fffff007f7fff80ffffffc07fffff81fff77fd1f7ff3f80ffbf07007d1e0000380c00000000e9006005ff0075dfff007ff7f70177ffff81ffffff01ffffff01ffffff01fff";
 when "00101110101" => data <= 768x"fffffffffffffffffffeffff7f70177ffff803fffff005fffff007fffff017f7fff00ffffff01ffffff81fff77f47f7fe3f00fffc1f007c7800007831010000139300800dff00554fff00ffc7f71177ffff03ffffff01ffffff01ffffff01fff";
 when "00101110110" => data <= 768x"ffffffffffffffffffffffff7f7d577ffff803fffff007fffff803fffff017f7fff00ffffff01ffffff81fff7ffc5f7feff03fffc7f00fdf80e00f8f00100507203000037d700551fff00ff8ff7117f7fff03ffffff01ffffff03ffffff01fff";
 when "00101110111" => data <= 768x"ffffffffffffffffffffffff7f7d777ffff817fffff007fffff003fffff017f7ffe00ffffff01ffffff01fff7f741f7fdff83fffc7f01fdf83e00f8f000005170020000755700045fff00fe1ff7107f5fff03ffffff01ffffff03ffffff017ff";
 when "00101111000" => data <= 768x"ffffffffffffffffffffffff7f7d777ffff817fffff007fffff003fffff007f7ffe00ffffff01ffffff01fff7f745f7f9ff83fff47f01fdf03e00f0f001004072020000775700447fff00fe17ff007f5fff03ffffff01ffffff03ffffff017ff";
 when "00101111001" => data <= 768x"ffffffffffffffffffffffff7f75177ffff807fffff007fffff003fffff007f7fff00ffffff01ffffff01fffdf7c7f7f8ff03fff07f01f5f03e00e0f0010000720200003f5f01551fff00ff07ff0577ffff03ffffff01ffffff03ffffff017ff";
 when "00101111010" => data <= 768x"ffffffffffffffffffffffff7f75177ffff807fffff007fffff003fffff007f7fff00ffffff01ffffff01fffdffc7f7f8ff03fff07f01f5f03e00e0f0010000720200003f5f01551ffe00ff07f70577ffff03ffffff01ffffff03ffffff01fff";
 when "00101111011" => data <= 768x"ffffffffffffffffffffffff7f7d7f7ffff83ffffff007fffff003fffff007f7ffe00ffffff01ffffff01fffff741f7f8ff83fff47f01fdf03e00f0f014004072020000374701451ffe00ff07ff057f7fff03ffffff01ffffff03ffffff017ff";
 when "00101111100" => data <= 768x"ffffffffffffffffffffffff7f7d7f7ffff817fffff007fffff003fffff007f7ffe00ffffff01ffffff01fff77f55f7feff83fffc5f01fdf01e00e0f100000073020000375701551ffe00ff87f7017fffff83ffffff01ffffff81ffffff01fff";
 when "00101111101" => data <= 768x"ffffffffffffffffffffffff7f7d177ffff803fffff007fffff807fffff007f7fff00ffffff01ffffff80fff77fd7f7fe3f01fefc1f007c780e00603101000013a300000ff700df8fff00ffffff0177ffff81ffffff01ffffff80ffffff017ff";
 when "00101111110" => data <= 768x"ffffffffffffffffffffffff7f7d177ffff803fffff007fffff807fffff017f7ffe00ffffff01ffffff80fff777d5f7ff3f81fffc1f007c780e007031000000138000000fd7005ddfff00fff7f70077ffff81ffffffc1ffffff80ffffff017ff";
 when "00101111111" => data <= 768x"ffffffffffffffffffffffff7f7f777ffff827fffff007fffff007fffff017f7ffe00ffffff01ffffff80fff7f741f7ffbfe3ffff1f007d7e0f007830010010108000000dd500454fff00fff7f70077ffff80ffffffc1ffffff80ffffff817ff";
 when "00110000000" => data <= 768x"ffffffffffffffffffffffff7f7f777ffff827fffff007fffff007fffff017f7fff00ffffff01ffffff80fff7f751f7ffbfe3ffff1f407d7e0700783c0100101020000005f50055cfff00fff7ff0077ffff80ffffffc1ffffff80ffffffc07ff";
 when "00110000001" => data <= 768x"ffffffffffffffffffffffff7f7d577ffff807fffff007fffff807fffff017fffff00ffffff01ffffff80fff7f751f7ffbfe3ff3f07007c1e0300681401000010a0006005f50075dfff80ffffff007fffff80ffffffc1ffffff80ffffffc07ff";
 when "00110000010" => data <= 768x"ffffffffffffffffffffffff7f7d177ffff803fffff005fffff807fffff007fffff00ffffff40ffffff80fff7ffd1f7ff9fe0ff3f07007c1e0300000400004000a00072edfd007fffff807ffff70077ffffc0ffffffc0ffffff80ffffffc07ff";
 when "00110000011" => data <= 768x"ffffffffffffffffffffffff7f7d177ffff803fffff001fffff803fffff007fffff00ffffffc07fffff80fff7ffd1f7ff9fe0ff3f07407c1e0380000400004000a00072edfd007fffff807ffff70077ffffc0ffffffc0ffffff80ffffffc07ff";
 when "00110000100" => data <= 768x"ffffffffffffffffffffffff7f7f777ffff803fffffc01fffff803fffff007fffff007fffff007fffff80ffffffc177ffdfe3ffbf47c07f1f03807c0c01000008200020057500757fff807ff7ff0077ffff80ffffffc1ffffff80ffffffc17ff";
 when "00110000101" => data <= 768x"ffffffffffffffffffffffff7f7d557ffff803fffffc01fffff801fffff001fffff007fffff407fffff80fff7ffd177ff8fe3ffff07417f5e03807e040100500a6000000ffd00715fff00fff7f70077ffff00ffffffc1ffffff80ffffff017ff";
 when "00110000110" => data <= 768x"ffffffffffffffffffffffff7f7d15fffff800fffff0007ffff800fffff005f7fff007fffff407fffff807ff7df5177ff8fe3ffff07017fde03007f8c4101550fe000000ffc00400ffe00f227f600777ffe00ffffff01ffffff01ffffff01fff";
 when "00110000111" => data <= 768x"fffffffffffffffffffebeff7f7c047ffff8007ffff0007ffff000fffff0057ffff007fffffc07fffff807fffdf5177ff8fe3ffff0701fffe02007fef50007f0ff000000ffc00400ffc00e007fc01755ffc00fffffd01fffffe03ffffff01fff";
 when "00110001000" => data <= 768x"ffffffffffff5ffffffc0c7f7f7c007ffff8003ffff0005fffe0007fff70057ffff803fffffc07fffff807ff7f7d077ffe3e3ffffc101ffff80007fef5000770fe0002a0ff000400ff800e007fc01711ffc01fbbffd01fffffe03ffffff03ff7";
 when "00110001001" => data <= 768x"ffffbffffffc041ffffc003f7f7c011ffff8001fffd0005fffe0023ffff00377fff803fffffc01ffffec03ff7fc717ffff860fffffc407fffe0003fff41007fdfc000330fd000400ff800e007fc01700ffe01fe8fff01ffdfff01ffffff01fff";
 when "00110001010" => data <= 768x"fffe003ffffc001ffffc000f7f7c001ffff8003fffc0017ffff801fffffc01fffffe00fffffc01fffffe03ff7ff7077ffffe07fffffc05fffc0803fff40001fffc0000bafd400500ffe007807ff017c0fff00fe2fffc1ff7fff80ffff7f017f7";
 when "00110001011" => data <= 768x"ffffa01fffff001ffffe001f7f7f001ffffe003ffff4007ffff800fffff4007fffff003fffff007fffff80ff7f7f41ffffff83ffffdf01fffe0e01fff50101f7fe00003fff500104fff003807f7107c0fffa07f0fffc07f5fffe07fff7fc07ff";
 when "00110001100" => data <= 768x"fffff83fffffd01fffff803f7f7f001fffff803fffff001ffffe003ffffd101fffff001fffffc01fffffc01f7f7f515ffffff0cfff5fc1c7ff07c087f7014017ff81803fffd00015fff801c07f7c01f0fffe03f0ffff01f0ffff83fdf7ff01ff";
 when "00110001101" => data <= 768x"fffffe1ffffff41fffffe01f7f7fc017ffff800fffffc01fffff801fffff001fffff800fffffc01fffffe01f7fff7417fffff8f3ffdff071ff83e060f701c045ff80c00fffdc4017fffc00807ffc01f0fffe01f0ffff01fcffff81fcfff7c1fd";
 when "00110001110" => data <= 768x"ffffff03fffffc07fffff0077f7f7005ffffe003ffffc007ffff8007ffff0007ffffe003fffff005fffff0037fff7115fffffe38ff57fc7cff83f838ff41f011ffc0e013fffc4007fffc00037ffc0151fffe0078ffff007cffffa0fcffffc07f";
 when "00110001111" => data <= 768x"ffffff80fffffc00fffff8007f7f7001fffff000fffff001ffff8000fff75001ffffe001fffff001fffff8007f7f7c01fffffe02ff57ff17ff01fe0eff017014ff80f00efffc5004fffc00007f7c0001fffe0000ffff001cffff803efffff03f";
 when "00110010000" => data <= 768x"ffffffa0fffffd00fffffc007f7f7c00fffff800ffffd000ffffc000ffffc000fffff000fffff400fffffc007fff7c00ffbffe00fe05ffc5fe01ff87ff01fd07ffb07802fff07007fff800027f7c0000fffe0000ffff0000ffff880efffff01f";
 when "00110010001" => data <= 768x"ffffffe0ffffff00fffffe007f7f7c00fffff800ffffd000ffffc000ffffd000fffff000fffffc00fffffc007f7f7c00fe0ffe00fc01ff41ff01ff87ff117d07fff07806fff05007fff800027f7c0000fffe0000ffff0000fffff80efffff01f";
 when "00110010010" => data <= 768x"fffffff8ffffff40fffffe007f7f7c00fffff800ffffd000ffffc000fffff000fffff800fffffc00fffffc007f5f7c00fe0ffe00fc01ff41fe01ff83ff117d07fff07006fff05007fff800027f7c0000fffe0000ffff5000fffff80cfffff01f";
 when "00110010011" => data <= 768x"fffffff8ffffff40fffffe007f7ffc00fffff800ffffd000ffffe000fffff000fffff800fffffc00fffffc007d5f7c00fc03fe00fc01ff40fe01ff82ff517d07fff07006fff05007fff800027f7c0000fffe0000ffff5000fffff808fffff01f";
 when "00110010100" => data <= 768x"fffffffeffffff40fffffe007f7f7e01fffff800ffffc000ffffe000ffff7000fffff800fffffc00fffffc007d177c00fc03fe00fc01ffc0fe01ff82ff507d07fff07006fff84007fffc00027f7c0000ffff0000fffff000fffff80cfffff01f";
 when "00110010101" => data <= 768x"ffffffe0ffffff00fffffe007f7f7500fffff000fffff000fffff800fffffc00fffffc00fffffc00fefffe007c177f00fc03ff80fc01ffc1fe00fe03ff707407fff82002fffc0007fffe00027f7f1001fffff800fffffc04fffff80efffff01f";
 when "00110010110" => data <= 768x"ffffff80fffffd00fffff8007f7f7000fffff800fffffc00fffffe00fff7f700fffffe00ff5fff00fe0fff807c077f50fc01ffe0fc007f41fe803c01f7f01001fffc0001fffd0000ffff80007f7fd400fffffc02fffffc07fffffc07fffff407";
 when "00110010111" => data <= 768x"ffffff00ffffff00ffffff807f7f7fc0ffffffe0ffffffc0ffffffe0f75ff7f0ff83fff0fc01fffcf8007ffe7d003f70fe000f80fe040700ff0e0000f71f0000ffbfe000ffffd000fffffb807f7f7fc1ffffff80ffffffc0ffffff80ffffffc0";
 when "00110011000" => data <= 768x"ffffffffffffffffffffffff7f57f77fffe3fffffd405ffffc000ffffc0007f7fe0003ffff40007cffc000387f714010fffff000fffff400ffebfe00ff01ff00ff83ffbeffc7fffcffc3fffc7f577f7cfffffffefffffffcfffffffcfffffffc";
 when "00110011001" => data <= 768x"ff0003ffff00007fff80003f7f400017ffe00003fffc0001fff80000fff01000fff83800fffffc00ffffff807f7f7fd0fffffffffffffffffffffffffffffff7ffffffffffffffffffeaffff7f007f7fff807fffffc0ffffffe1fffffff1ffff";
 when "00110011010" => data <= 768x"ffff0030fffc0014fff000027f741401ffffbe00ffffff40ffffffe0fff7fff5ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7fffebffffff007fffff007fffff0077ff";
 when "00110011011" => data <= 768x"fffffffafffffffdffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ff77f7fff803fffff007fffff803fffff407fff";
 when "00110011100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffbbfffff801fffff801fff7fc01f7fffe03ffffff07fffffe0fffffff17fff";
 when "00110011101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f75577fffc00fffffc00fffffc00fffffd01ffffff03ffffff07ffffff83fff7f757f7fffffffffffffffffffffffffffffffff";
 when "00110011110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff017ffffe007ffffc007ffffe00fff7f701f7ffff83ffffff87ffffff83ffffffd77ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110011111" => data <= 768x"ffffffffffffffffffffffff7f777f7ffff03fffffc007ffffe003fffff007fffff00ffffff01ffffff83fff7f743f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100000" => data <= 768x"fffffffffff57fffffe00fff7f70077fffe007fffff007fffff00ffffff01ffffff83ffffffc7fffffffffff7f7fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100001" => data <= 768x"fff0bffffff01fffffe003ff7f71057ffff00bfffff007fffff83ffffff07ffffffa7fffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100010" => data <= 768x"ffe03fffffe01fffffe003ff7ff0057ffff00bfffff017fffff83ffffff077ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100011" => data <= 768x"fff3ffffffc05fffffe00fff7f7005fffff003fffff005fffff80bfffff057fffff83fffffff7fffffffffff7f7fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100100" => data <= 768x"ffffffffffffffffffffffff7f75ffffffe03fffffc017ffffe003fffff005fffff007fffff015fffff03fff7f757f7ffffffffffffffffffffffffffff7ffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffffffe3ffffffc05fffffe007ff7f7001fffff003fffff005fffff00ffffff07ffffffe7fffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "00110100110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffffffffffffffff7f7fff7ffffbffffffc17fffffe03fffff7017ffffe003fffff005fffff005ff7f70157ffff03ffffff47ffffffefffffff7f7ff";
 when "00110100111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080000003d4000003ff000001dfc00003ffe00001f7f00000ffe80001ffd00001fea00001fc000";
 when "00110101000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000788000007dd000003ef0000077f400003fee00001fdf40000fff00001fff40001fea80001f4000";
 when "00110101001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fec000007470000062f80000777400003b8700001ff700001fff80001fff40001fe380001f4000";
 when "00110101010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000008000000100000001000000050400000e060000140740000c278000051514000798380001df740001fffe0001dff40001ffbc000171000";
 when "00110101011" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000400000004000000040000000e00000004040000000600001017c0000813800005101400078e380001df741003effe0001d7fd0001ff8a000171040";
 when "00110101100" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000180000001400000002000000000000000000000000040000200380001001c000180800001d0c14000f8f380001c7740003effe0001f7d70001fbca000171040";
 when "00110101101" => data <= 768x"000000000000000000000000000000000300000007c00000038000000300000003000000010000000000000000000000000000000400100000001800070054000380400001d045d000f87180003c7340003ef7e0001d7d70001fbca000171450";
 when "00110101110" => data <= 768x"000000000000000000000000140000001e00000007000000030000000100000000000000000000000000000000000000000000000000100008000c00050000000380200001d0715000f87080007c71c0003e73e0001d7d70001fbcb000151450";
 when "00110101111" => data <= 768x"0000000000000000000000005500000038000000000000000000000000000000000000000000000000000000000000000000000000001c0008000c00150010010f80106007d0505000f87080007c71c000383be0001f3d70001fbcb000151450";
 when "00110110000" => data <= 768x"000000000400000000000000140000003800000010000000000000000000000000000000000000000000000000000000000000000000000000000c0004000500060000000740045403f0383e017c3c50003e3ce0001d1df0000f8ef80017df1c";
 when "00110110001" => data <= 768x"0000000000000000000000000500000002000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000001c000000000005000000048000000750544003f87cf001fc755";
 when "00110110010" => data <= 768x"000000000000000000000000000000000020000000f0000000f0000001d0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000008000000040000000000010000";
 when "00110110011" => data <= 768x"00000000000000000000000000000000000000000010000000380000001c000000380000001c00000008000000050000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
 when "00110110100" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000140000000e000000074000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110110101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000004000000380000007000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110110110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000100000000800000010000000080000001c00000018000000100000000000000000000000000000000000000000000000000000000000000000000";
 when "00110110111" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000740000003e0000000600000004000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111000" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000020000000f0000001e000000170000003e0000007400000060000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000010000000380000007c0000003c0000003c000000380000001c00000008000000040000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111010" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000150000000f80000007c0000007e0000005500000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000010000003b00000075000000fc000001fc00000020000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111100" => data <= 768x"0000000000000000000000000000000000000000000000000000000000004000000080000000c0000003c0000001c0000003c0000007c00000038000000300000002000000000000000000000000000000000000000000000000000000000000";
 when "00110111101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000080000000500000003c0000003c0000003e0000001c0000000c000000060000000200000000000000000000000000000000000000000000000000000000000";
 when "00110111110" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000001c0000003e000001770000033f8000001440000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00110111111" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000018000001d0000003e0000007c000000780000007c00000068000000400000008000000000000000000000000000000000000000000000000000000000000";
 when "00111000000" => data <= 768x"00000000000000000000000000000000000000000001000000018000000100000001000000050000000780000007c0000007e0000007c00000038000001040000000400000004000000000000000000000000000000000000000000000000000";
 when "00111000001" => data <= 768x"00000000000000000000000000000000000000000000000000000000001000000030000000140000000fc000000740000007fa000007d5000003c000000100000000000000000000000000000000000000000000000000000000000000000000";
 when "00111000010" => data <= 768x"000000000000000000000000000000000000000000000000000008000000140000001000000150000003e0000007f1000007e000001fc0000063c000004100000000000000000000000000000000000000000000000000000000000000000000";
 when "00111000011" => data <= 768x"0000000000000000000000000000000000020000000100000001000000010000000100000001c0000003e0000007f0000003e0000001f0000001e000000140000001000000010000000300000001000000000000000000000000000000000000";
 when "00111000100" => data <= 768x"0000000000000000000000000000000000000000000000000000000000010000006000000055c000000fe000000770000003f0000005f0000000a000000010000000080000000400000000000000000000000000000000000000000000000000";
 when "00111000101" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000180000005c1000007ff000007f5000007e000001fc00000310000004100000000000000000000000000000000000000000000000000000000000000000000";
 when "00111000110" => data <= 768x"00000000000000000000000000001000000030000000500000006000000040000003c0000007c000000fe0000007c000000fc0000007c0000007a000001100000001000000010000000180000001000000000000000000000000000000000000";
 when "00111000111" => data <= 768x"000000000000000000200000007100000038000000140000000c00000007d0000003e0000007c000000fe000001ff000001ff000001ffc00000fee000017d7400003838000010140000000000000000000000000000000000000000000000000";
 when "00111001000" => data <= 768x"000000000000000000000000000140000003c0000007c0000007e00000075550001ffff0017fd5500bffe00017077000080ff800001ff400003ff800003ffc00003ff800001ff000000fe0000007400000010000000000000000000000000000";
 when "00111001001" => data <= 768x"0000000000014000000fc000001f4000000fc000000fc000000fe000000575400003ff000007f000001fe000001f7000003be0000015f000003fe0000077740000e7fe0001c7fc00038ffe00071f7d00023ffe00041ffc00001ffc000007f000";
 when "00111001010" => data <= 768x"00000000000000000000000000074000000fc0000007c000000fc0000007c0000007c0000005c0000003e000000750000007f8000007f4000007e000000760000007e000001fc000000fe000001ff0000027f8000047fc000007fc0000177400";
 when "00111001011" => data <= 768x"000000000000000000000000000000000000000000054000000780000007c000000780000007c0000007800000070000000380000007c0000007e0000007c0000003e0000007c0000007e000000770000007f0000007d0000013e0000037c000";
 when "00111001100" => data <= 768x"000000000000000000000000000000000000000000000000000380000007c000000780000007c0000007c00000074000000380000007c0000003c0000003c0000003e0000001f0000003f80000075c000007e8000007c4000007e0000017c000";
 when "00111001101" => data <= 768x"000000000000000000000000000000000000000000000000000380000007c000000780000007c0000007c00000074000000380000007c0000003c0000001c0000003f0000001f4000007e800000744000007e0000007c0000007e0000007f000";
 when "00111001110" => data <= 768x"000000000000000000000000000000000000000000000000000380000007c000000780000007c000000fc00000074000000380000007c0000003e0000001f0000001f8000001dc000007e800000760000007e0000007c000000fe0000007f000";
 when "00111001111" => data <= 768x"000000000000000000000000000000000000000000000000000380000007c000000780000007c0000007c00000070000000380000007d0000003f0000001f0000001f0000005f000000fe0000007f0000007f0000007d000000fe0000007f000";
 when "00111010000" => data <= 768x"000000000000000000000000000000000000000000000000000380000007c000000780000007c0000007c00000070000000f8000000fc0000007e000000170000003f0000005f000000ff800001750000007e0000007e000000fe0000017f000";
 when "00111010001" => data <= 768x"000000000000000000000000000000000000000000000000000280000007c0000007c0000007c0000007c00000074000003fe000001ff000000bf0000003f0000003f8000005f000000fe000001741000007e0000007c000000fe0000017f000";
 when "00111010010" => data <= 768x"000000000000000000000000000000000000000000000000000080000007c0000003e0000007c0000003e0000011c000003fe000007ff000000ff0000007f0000003e0000007d0000007f000000770000007e0000007c000000fe0000017f000";
 when "00111010011" => data <= 768x"000000000000000000000000000000000000000000000000000080000003c0000003e0000001f0000003e0000001c000001fe000001ff000002fe0000007c0000003c0000017c0000007f000000770000007e0000007c000000fe000001ff000";
 when "00111010100" => data <= 768x"0000000000000000000000000001000000000000000100000003e0000001f0000003e0000001f0000001e00000014000000fe000001fe000001fc0000017c000003f80000007c0000007e00000077000000fe0000007c000000fe000001ff000";
 when "00111010101" => data <= 768x"0000000000000000000000000000000000000000000140000001e0000001f0000003e0000001f0000000e0000005c000000fe000001fc000003fc0000057c000000380000007c0000007f0000007f000000fe000000fc000000fe000001ff000";
 when "00111010110" => data <= 768x"00000000000000000000000000000000000000000001c0000003e0000001f0000003e0000001f0000000e00000174000007fc000015fc000000f800000078000000380000007c0000007e00000077000000fe000001fc000000fe000001ff000";
 when "00111010111" => data <= 768x"00000000000000000000000000000000000080000001c0000003e0000001f0000003e0000041f00000e3e0000177c000000fc0000007c000000f800000070000000780000007c0000007e00000077000000fe000000fc000000fe0000017f000";
 when "00111011000" => data <= 768x"00000000000000000000000000000000000080000001c0000003e0000001f0000283e00005f5f00000bfe0000017c000000fc000000fc000000f800000070000000780000007c0000007e00000077000000fe0000007c000000fe0000017f000";
 when "00111011001" => data <= 768x"00000000000000000000000000010000000080000001c0000001e0000141700000e1f0000075f000000fe0000007c000000fc000001fc0000007800000070000000780000007c0000007e000000770000007e0000007c000000fe0000007f000";
 when "00111011010" => data <= 768x"0000000000000000000000000001000000000000000140000081e0000051f0000031f000001df000000fe00000074000001fc0000017c0000007800000070000000780000007c0000007e000000770000007e0000007c0000007e00000077000";
 when "00111011011" => data <= 768x"00000000000000000000000000000000000000000040400000c1e0000071f0000039f000001df000000fe00000174000001fc0000017c0000007800000070000000780000007c0000007e000000770000007e0000007d0000007e0000007f000";
 when "00111011100" => data <= 768x"0000000000000000000000000000000000000000004140000061e0000071f0000039f000001df000000fe000001f4000001fc0000017c0000007800000070000000780000007c0000007e0000007f0000007e0000007d0000007e0000007f000";
 when "00111011101" => data <= 768x"00000000000000000000000000000000000000000041c0000061e0000071f0000039f000001df000000fe000001fc000001fc0000017c0000007800000070000000780000007c0000007e0000007f0000007e0000007d0000007e0000007f000";
 when "00111011110" => data <= 768x"00000000000000000000000000000000000000000041c0000021e0000071f0000031f000001df000000fe0000017c000000fc000001fc0000007800000070000000780000007c0000007e0000007f0000007e0000007e0000007e00000077000";
 when "00111011111" => data <= 768x"00000000000000000000000000010000000180000001c0000003e0000017f0000033f0000071f000003ae00000174000000fc000001fc000001f80000017c000000780000007c0000007e000000770000007e0000007e000000fe00000077000";
 when "00111100000" => data <= 768x"00000000000000000000000000010000000380000007c0000007e0000007f0000003e0000007f0000003e00000175000001ff000001ff000001ff0000017d0000007c0000007c0000007e000000770000007f8000007f000000ff000001ff000";
 when "00111100001" => data <= 768x"00000000000000000000000000170000000fe000001fc000000fe000001ff000000ff0000007f0000003e00000075000000ff800001ffc00001ffc00001ffc00001ff800001ffc00000ff800000770000007fc000007fc00000ffc00001ff400";
 when "00111100010" => data <= 768x"000000000000000000000000001f4000001fe000001ff000001ff0000017f000001ff0000007f0000007e0000005d000000ff800001ffc00000ffe00001ffc00000ff8000007fc000003f8000017fc00000ffc000007fc000007fe000007fc00";
 when "00111100011" => data <= 768x"000000000000000000000000001f4000001fe000001ff000001ff0000017f000001ff0000017f0000007f0000007d1000003f3800007ffc0000fff800007ff000007fc000007fc000003fe0000017f00001bff00001fff00000ffe000007f400";
 when "00111100100" => data <= 768x"00000000000001000000000000174100000ff100000ff100000ff980001ff100000ff9800007fdc00003f8c0000171c00003fb800007fdc00003ff800003f7000003fe000001fc000001ff000001ff000009ff80001fff00000ffe000007fc00";
 when "00111100101" => data <= 768x"000000000000004000000080000750400003f8000007fc400003fc400007fc400003fe600005fc700000fe60000174700000fee00001ffc00001ffc00001ffc00000ff8000007f000000ff8000007fc000027fe00007ffc00003ff8000017f00";
 when "00111100110" => data <= 768x"0000000000000040000000200001f4010001fe200001ff100001ff200001ff100001ff3800017f1000007f3800005f1000003f3800007f7000007fe000007ff000007fe000007fc000003fe000001f7000033ff00001fff00001ffe000017f40";
 when "00111100111" => data <= 768x"000000000000001000002000000175100000ff1000007f100000ff980001f7900000ff9800007fdc00003f8c0000171c00003f9800007fdc00003ff800003ff000003fe000001fc000001fe000001f700000bff80001fff00000ffe000007fc0";
 when "00111101000" => data <= 768x"00000000000000100000200000007f100000ff0000007f140000ff8800017fdc0000ff8c00007fdc00003f8e0000171c00003f9c00005fdc00003ff800001ff000003ff000001fd000001fe000001f700000bff80001fff00000ffe000007fc0";
 when "00111101001" => data <= 768x"00000000000000000000380800007f000000ff8000007fc40000ff8c00007fc400007fce00005fcf00003f8e0000175700003fde00001fdc00003ff800001ff000001ff000001ff000000fe000011f700000fff80001fff00000ffe000007fc0";
 when "00111101010" => data <= 768x"000000000000100400003e000000770400007f8000007fc400007fc600007fc700003fe700001fc700001f870000174700001fef00001fdc00001ffc00001ff000001ff000001ff000000fe000011f700000fff80001fff000007fe000007fc0";
 when "00111101011" => data <= 768x"000000000000540400003f8000007fc400003fc600007fc400007fe200007f7700003fe300001fc700000f8700001f4700001fee00001fdc00000ffc00001ff000000ff000001ff000000fe000015f700000fff800007ff000007fe000007fc0";
 when "00111101100" => data <= 768x"0000000000000000000000000000000000000000000570000007f8000007fc000007ff000007ff000007fe00000575000000f800fd547c000ffefe000177f7c0003fffc00005ffc40000fffe00007f7f00003fbe00007fdc00003ff800007f70";
 when "00111101101" => data <= 768x"0000000000000000000000000000010000000000000000000000bc000001ff000001ff000001ff540001fffe00017f7400007fe000007fc000002f80000007c000000fc000001fc000000fe00000177000000ff8000007fd000003ff000001ff";
 when "00111101110" => data <= 768x"00000000000000000000000000000000000000000000000000000007000000170000001f0000005f0000003f0000001f0000000f0000001f0000000f000000150000000000000001000000000000000100000000000000000000000000000000";
 when "00111101111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005400000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000554000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000057400000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015500000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000232000005550000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110100" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100003fff00005555000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000040000000c0005555d0003ffff0000041c0000000c000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110110" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000577f00000bff0000000500000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00111110111" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000020001577f0003ffff0000455700000003000000070000000f0000001f0000000f0000001f0000001f0000001f0000000f00000017";
 when "00111111000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f0001577f03ffffff0555f55c0000e03c0001707d0001f87e0001f47d0003f8ff0001747f0003f87e0001f47d0001f83e0001f07d";
 when "00111111001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000001000000070000005d000003ff01015ff303bffbe37ffdd1d701c0c1e301c1d1f303e3e3f307d1f1f103e3e1e103f1715103e1e1e101c1d1c101e1e0c001c1d1c0";
 when "00111111010" => data <= 768x"00000000000000000000000000000000000000000000000100000000000001c0000003e000001f700000fe380017f71d03ff8f3effd1c77fe0c3cfff71d3c775f1e3c73bf1f1c717f1e3c63b71d1c717f0e1821371c1401160c1800370411001";
 when "00111111011" => data <= 768x"0000000f000000070000000f000000070000000f0000001f0000003f0000005f0000e03b0001f01d000f3818015f1c1c0bf39e08fd47df01b8e3bf8311731dd738f3bbbf7c711ddf38e11bbf1461117f386003bf1040011f1800019f10000117";
 when "00111111100" => data <= 768x"0000003f000001ff000003ff0000017f000003ff000001ff000003ff000007f7000003ff001c077f007e072f05f707173f33823fd477407f8e7760ffd777757f8e2377ffc477747f8e226eff0411777f840026ff040045ff000026ff000005ff";
 when "00111111101" => data <= 768x"00000020000015f400001ffc00001f7c00003ffc00001ffc00001ffe0000177400003ffe004077f401e033f0177171713f3833f8771407fc23be0ffe733357f773337fff711747ff2026efff3117777f20026fff000447ff00000ffe000017ff";
 when "00111111110" => data <= 768x"000000000000054000001fc000007f600000ffe00001ffc00000ffe000007ff00000ffe00001dfc00300cf801541c700f8e08fe0ccd01ff08cd83ff0d5dd77f5cc9bbffbc45d1ff1809bbffb00113f71001b3ff900117ff100003ff0000077f0";
 when "00111111111" => data <= 768x"000000000000040000003f8000017fc00003ff800001ffc00001ffc00001f7c00001bfc000015f400e03bf0017011700f9811f805d417fc099a07fc011157ff599b2ffe611767ff780367fe601377f7700227fe200047fc40000ffe0000077c0";
 when "01000000000" => data <= 768x"000000000000040000003f8000017f000003ff800001ffc00003ff800001ffc00003bfc000017f400e03bf0017011700f9833f005d417fc09ba07fc011157ff59932ffe611747fe400367fe601367f6400227fe600047fc40000ffe000007fc0";
 when "01000000001" => data <= 768x"000000000000040000003f8000017f000003ff800001ffc00003ff80000177c00003ffc000017f400e03bf0017011700f9833f0059417fc09ba07fc0111577f59932ffe611747fe500367fe601367f6400227fe600047fc40000ffe000007fc0";
 when "01000000010" => data <= 768x"000000000000000000003f0000017f000003ff800003ffc00003ff80000177c00003ff8000017f400e03be0017011700f9833f8059417fc09ba07fc0111577d59932ffe611747fc500267fe601367f4400227fe600047fc40000ffc0000077c0";
 when "01000000011" => data <= 768x"000000000000000000003f0000017f000003ff800007ffc00003ff8000017fc00003ff8000017f400e03be0017031700f1833f0059417fc09ba07fc0111577d59932ffe411747fc50026ffee01347f4400267fe400047fc40000ffc0000077c0";
 when "01000000100" => data <= 768x"000000000000000000003e0000017f000003ff800007ff000003ff8000017fc00003ff8000017f400e03be0017031700f1833f0059417fc09ba07fc0113577d59936ffe411747fc50026ffec01347f450026ffc400047fc40000ffc0000077c0";
 when "01000000101" => data <= 768x"000000000000000000003e0000017f000003ff000007ff000001ff8000017f000003ff0004077f000e033e0011031d00f9833f005d407fc099a07fc0d1157f558932ffe511767fc580267fec00147f450022ffc000047fc40000ffc0000177c0";
 when "01000000110" => data <= 768x"00000000000054000000fe000001ff000003ff000001ff000003ffc00007ffc00003ff0001057d000f033e005d431d00ece03f004dd07fc0cd987fcbd5957fd589b2ffefc1177fc580367fec00177f450002ffc000047fc40000ffc00001ffc0";
 when "01000000111" => data <= 768x"000000000000140000007e0000007f000000ff800001ff000003ff800001ffc00001ff800101ff000e81be007441150026e03f0044d07fc06cc87fef45d57f55409b7fef44177fc500127fec00177f450002ffc000007fc00000ff800001ffc0";
 when "01000001000" => data <= 768x"0000000000001c0000007f0000017f000001ff800001ff000001ff8000017fc00000ff8001007f000ec03e007740550026703f0077507f0126ccffff745d7f55201b7fef40597fc5001bffec00137f450002ff8000017fc00000ff800001ffc0";
 when "01000001001" => data <= 768x"0000000000001c0000007f0000017f000001ff800001ff000001ff8000017fc000007f8001007f000ec03e0077401d0022703f0077507f0532ecffff365d7755225bffed005d7fc5000bffec00117f450003ff8000017fc00000ff800001f700";
 when "01000001010" => data <= 768x"0000000000005c0000007f0000017f000001ff800001ff000003ff800001ffc000007f8001007f000e803e0074401f0026603f0077507f052268ffff335d7f55223bffed105d7fc5000bffec00117f450001ff800001ff800000ff800001ff00";
 when "01000001011" => data <= 768x"0000000000005c000000fe0000017f000001ff800001ff000003ff800005ff4000007f8001007f000e803e0074401d0066603f0077507f056268fffb315d7f5d303bffed105dff4d000bffc800057f450001ff800001ff000000ff800001ff00";
 when "01000001100" => data <= 768x"0000000000005c000000fe0000017f000001ff000001ff000003ff800005ff4000007f0005007f000e803c0074401d0066603f0067507f0562e8fffb735d7f5d323bffe9105dff4d000bffc800057f450001ff800001ff000000ff800001ff00";
 when "01000001101" => data <= 768x"00000000000054000000fe000001ff000001ff000001ff000003ff000005ff000000ff0005007d000c80380074401d0066e07f0046d07f1566c8fffb7657ffd3227bffdb105f7fd9000bffc800117f400001ff800001ff000000ff800001ff00";
 when "01000001110" => data <= 768x"00000000000050000001f8000001fc000003fe000007fc000007fe000007f7000001fc000501f4000d00700055417c01ada1fe0375d5fd55ecbfffad6575ff7520b6ff244015ff640026ff200015ff010001ff000001ff000003fe000007ff00";
 when "01000001111" => data <= 768x"00000000000140000003e00000077000000ff8000007f000000ff8000017f1000003f0000001c0040380e00e15c170131da3f27b5d17fd5de9b7ffe97177fd75e82ff9204045dd00000bec000103f5000007f8000007fc00000ffc000017fc00";
 when "01000010000" => data <= 768x"0000000000050000000fe000001f7000001ff000001fd000003fe000001fc0000007c0000005c100003b8380005f55c001fffe7001f7fd1c038fe80f171ff0013e07e0007007e000f007e0005007e000001fe0000017e0000027e0000077f000";
 when "01000010001" => data <= 768x"0000000000054000000fe000001f7000001ff000001fd000003fc0000017c000000fe0000007c4000007c20000075c000007fe000007fc00000ffe000007fd000007fe000007dc000007fc00000754000007fc000017fc00000ff8000017f000";
 when "01000010010" => data <= 768x"0000000000054000000ff000001ff000000ff800001ff400001ff0000017f000000ff0000145f00001c7e01803777075023ffbae0007f5050007e801000770010007e0000007f0000007e00000077000000fe0000007f000000ff0000017f000";
 when "01000010011" => data <= 768x"00000000000000000003e0000007fc00000ffc000007fc00000ff8000017f8000007f8000005dc003c03d80075077074c3fffbbf0147f7d5000fe0010007f0000007f0000007f000000ff00000077000000fe000001ff000000ff000001ff000";
 when "01000010100" => data <= 768x"00000000000000000002c0000007f0000007fc000007fc00000ffc000017f4000007ec000005cc0008018c0015077010fbbff03cc747f7d5800ff3830007f001000ff0000007f000000ff000001f7000000ff000001ff000001ff0000017f000";
 when "01000010101" => data <= 768x"0000000000000000000280000007f0000007f8000007fc00000ffc000017f4000007ec000005c400000384001507f0502d2ff0f855dff754838ff3870517f111000ff000000ff000000ff000001f7100001ff8000017f000001ff8000017f000";
 when "01000010110" => data <= 768x"0000000000000000000280000007f0000007f8000007fc00000ffc000017f4000007e8000005cc0000038c001407c050672fe0f8755ff55485cff70f1157f117800ff000001ff000001ff000001750000037f8000077f000006ff800005ff400";
 when "01000010111" => data <= 768x"0000000000000000000280000007d000000ff8000007fc00000ff8000017fc000007f8000005dc000003880014074050262fe0f8555ff5f59befef0f515ff417403ff003401ff00003b7f00001f750000087f8000007fc00000fe800001ff400";
 when "01000011000" => data <= 768x"0000000000000000000280000007d000000ff8000007fc00000ff8000017f8000007f8000005dc00000388001407c050272fe3fa55dffd559abfff2c415ff411201ff0020117f00403e7f000014750010007f8000007fc00000ff800001ff400";
 when "01000011001" => data <= 768x"0000000000000000000380000007d000000ff8000007fc00000ff8000017d0000007f8000005dc00000388001407d154262ffbfa55dfdd55cabffaa6415ff405200ff0010017f0018033f00005c750000307f8000007fc00000ff8000017f400";
 when "01000011010" => data <= 768x"00000000000000000003c0000007f000000ff8000007fc00000ff8000017f8000007f8000005dc000003880014075154262ffb6a55dffd51dabffb4a505ff113200ff0020017f0000033f000014750000307f8000007fc00000ff8000017f400";
 when "01000011011" => data <= 768x"00000000000000000003c0000007f000000ff8000007fc00000ff8000017f8000007f8000005dc000003880014074054272ffb2e55dff54dd0bff92b501ff101000ff0010017f0000033f800014750010387f8000407fc00000ff8000017f400";
 when "01000011100" => data <= 768x"00000000000000000003c0000007f000000ff8000007fc00000ff8000017fc000007f8000005dc00000388001507f054272ffbae555ff53580bffda75117f511000ff0000017d0000033f800014771000387f8000407fc00000ff8000017f400";
 when "01000011101" => data <= 768x"00000000000000000003c00000077000000ff8000007fc00000ff8000017fc000003f8000005dc00080388001507f054272ff0ae555ff515a9afe4970117f511000ff0000017f0000033f800014750000387f8000407fc00000ff8000017f400";
 when "01000011110" => data <= 768x"00000000000000000003e0000007f000000ff8000007fc00000ff8000017fc000003ec000005cc00080388001507f050252ff02ed55ff515a9aff6970117f451000ff2000017f0400033f800014770000387f8000407fc00000ffc000017f400";
 when "01000011111" => data <= 768x"00000000000000000003e0000007f0000007f8000007fc00000ffc000017f4000003ec000005cc00080388001507701065aff024f55ff515a9aff6970157f455000ff2010017f0000033f80001475d000387ee000407f700000ff3000017f310";
 when "01000100000" => data <= 768x"00000000000000000003e0000007f0000007f8000007fc00000ffc000017f4000003ec000005cc0008038c001507601065aff024d55ff515a9aff6ad0157f515800ff2010017d0410033ec80014747000387e0000407f000000ff0000017f000";
 when "01000100001" => data <= 768x"00000000000000000003e0000007f0000007f8000007fc00000ffc00001774000003ec000005cc0008018c0015074010e7aff024d55ff535a5aff6ad1547f715800ff283001fd0010033ec80015747400387e0000507f000000ff0000017f000";
 when "01000100010" => data <= 768x"00000000000040000003e0000007f0000007fc000007fc00000ffc000017f4000003ec000005c40018018c0075074014b7aff024955ff575a5aff6a9d547f501800ff2020017d0000037ec00015747000387e1a00507f040000ff0000017f000";
 when "01000100011" => data <= 768x"00000000000140000007e0000007f0000007fc000007fc00000ffc000017f4000003ec000005c40018038c0075074014a7aff026955ff57595aff6a9d577f511802ff2024017d4040037ec00015747010387e1800507f050000ff0000017f000";
 when "01000100100" => data <= 768x"00000000000140000007e00000077400000ffc000007fc00000ffc000017f4000003ec000005c40018038c0075074014a72ff026155ff57595aff6a9d577f551802ff102401fd4040037ec00015747000387e3800507f050000ff0000017f000";
 when "01000100101" => data <= 768x"00000000000140000007e00000077400000ffc000007fc00000ffc000017f4000007ec000005c40000038c0054074014e72ff026155ff575b5affcadd577f50180aff103401fd5000037ec00015747000387e3800507f050000ff0000017f000";
 when "01000100110" => data <= 768x"00000000000140000007e00000077400000ffc000007fc00000ffc000017f4000007ec000005c40000038c00540744146f2ff026755ff555a5affcadd537f50580aff103401fd5010037ec00017747000387e3800507f050000ff0000017f000";
 when "01000100111" => data <= 768x"00000000000540000007e00000077400000ffc000007fc00000ffc000017f4000007ec000005cc0000038c00540744146e2ff036755ff515adaffcac9537f515802ff081401ff501003fec00017747000387e3800707f050000ff0000017f000";
 when "01000101000" => data <= 768x"00000000000540000007e0000007f400000ffc000007fc00000ffc000017f4000007ec000005cc0000038c00540744146a0ff0327d5ff515a92ffeb41577f595812ff481011ff401003fec00017747000387e3801707f050000ff000001ff000";
 when "01000101001" => data <= 768x"0000000000054000000fe00000077400000ffc000007fc00000ffc000017f4000007ec000005cc0000038c00140744146a0ff0325d5ff515292ffe964177f5d5a12ff480011ff400003fec00017767000387e3801707f050000ff000001ff000";
 when "01000101010" => data <= 768x"0000000000054000000fe0000007f400000ffc00001ffc00000ffc000017f4000007ec000005c40000018c00540740146a0ff0325d5ff5d56b6ffe964177f5d5012ff282011ff440003fec00007767010387e3801707f050080ff000001ff000";
 when "01000101011" => data <= 768x"0000000000054000000fe00000077c00000ffc00001ffc00001ffc000017f4000007ec000005c40000018c00540740146a0fe0325d5ff5576b6ff69651577755032ff282015ff440003ffc000077670003c7e3801707f1500c0ff020001ff000";
 when "01000101100" => data <= 768x"0000000000054000000fe00000077c00000ffc00001ffc00001ffc000017f4000007ec000005c40000018c005407c0144a0ff0325d5ff5576b6ffe9651577755026ff282015ff440003ffc000077670003c7e3801707f1500c0ff020001ff000";
 when "01000101101" => data <= 768x"000000000007c000000fe00000077c00000ffc00001ffc00001ffc000017f4000007ec000005c40000018c005007c0144a0ff0335d5ff5576b6ffede51577755026ff282415ff040003ffc000077770003c7e3801707f1500c0ff0200017f000";
 when "01000101110" => data <= 768x"000000000007c000000fe00000077c00000ffc00001ffc00001ffc000017f4000007ec000005c40000018c005007c014ca0ff0335d5ff5576b6ffad653577755025ff282415ff040003ff8000077770002c7e3801707f1400e0ff0200017f000";
 when "01000101111" => data <= 768x"000000000007c000000fe0000007fc00000ffc00001ffc00001ffc000017f4000007ee000005c400000184005007c015ca0ff0335d5ff5576b4ffad653577755025ff282415ff040003ff8000077770002e7e3800707f1400e0ff0200017f000";
 when "01000110000" => data <= 768x"000000000007c000000fe0000007fc00000ffc00001ffc00001ffc000017f4000007ee000005c400000384005007c015ca0ff0335d5ff5576b4ffad6535777550b5ff280415ff040003ff8000077770002e7e3801707f1c00e0ff0200017f000";
 when "01000110001" => data <= 768x"0000000000054000000fe00000077400000ffc00001ffc00001ffc000017f4000007ee000005c40000018c005007c514480fe0335d5ff5576b7ffa9e5357f7552b7ff280415ff455003ffc00057777412fe7e3e01d07f174000ff0000017f000";
 when "01000110010" => data <= 768x"0000000000054000000fe00000077400000ffe00001ffc00001ffc000017f400000fee005005c40478038e1a5d0744576bafef925d5ff4564b7ffed2515ff650025ff200005ff400003ff80015777f743fe7eff81547f150000ff0000017f000";
 when "01000110011" => data <= 768x"000200000007d0000007f00000077400000ffe00001fff00000ffe000007f4103807fe266405c555e9a38fb65d57d5d74b2ff692417ff450027ffa80015ff400001ff800001ffc00003ff80004777d152ee7ef3c5fc7f5fc0f0ff0f80017f000";
 when "01000110100" => data <= 768x"fffefffffffc1ffffff80fff7f70057fffe001fffff001fffff001fffff001f7eff809e3d5fc515912ee304817501145b680032f74c00175fc8003bffdd0057fffe007ffffc007ffffc803fff75011dfb31818cbc0501c01e8f00e03fff00777";
 when "01000110101" => data <= 768x"fffe3ffffffc1ffffff80fff7f70057fffe001fffff001fffff001fffff001f7eff809e3d5fc515912ee304817501145b680032f74c00177fe8003bff5d00777ffe007ffffc007ffffc803fff75011dfb31818cbc0501c01e8f00e03fff00777";
 when "01000110110" => data <= 768x"fffc3ffffffc07fffff807ff7f7005ffffe000fffff001fffff001fffff001f7e7f809e355fc515d12ec304815501145b680032f74c0017dfec003bff5d00777ffe007ffffc007ffffc803ff775011ffb31818ebc0501c01c0f00e03f5f00757";
 when "01000110111" => data <= 768x"fff80ffffff407fffff807ff7f70017fffe000fffff001fffff000fffff101f7e7f809eb15fc515d928c306815501145b480032dd5c0017dfec003fff7c00777ffe003ffffc007ffffc803ff771011f7b618086f44501c4180f00e01f5f00757";
 when "01000111000" => data <= 768x"fff807fffff007fffff800ff7f50017fffe000fffff001fffff008ffdff105f7a3f808e815dc5545a688302815501105b480032dd5c0017dfec003ffffc0077fffc003ffffc007ffffc003ff7f1011f76610086644501c4080f00e00d5f00755";
 when "01000111001" => data <= 768x"fff803fffff0057fffe000ff7f40007fffe000fffff0047ffff000ffd7f1057123fc08e6555c5445a48810a415100115b480012dd5c0017dfec003fff7c00777ffc003ffffc001ffff8003ffff1011f7ee10087744500c1400f00e0051f00741";
 when "01000111010" => data <= 768x"fff0027fffd0007fffc0007f7fc0007fffe0007ffff0047ffff004f957f5047563fe3822455c5014218000a435100115b98001afd5c0017dff8003fff7c003ffff8003ffffc001ffff8003ffff101177de30083b54500c1100f00e0001f00740";
 when "01000111011" => data <= 768x"ffe0003fffc0007fffc0003ffff0007fffe0027ffff0047d1ff8047857f414714bbe3812451450500980008261000115a90001bffd0001dfff8001fff7c001f7ff8003ffffd001ffff8001ff7f10117fbe30083d1470041d00e00e0001f00741";
 when "01000111100" => data <= 768x"ff80003fffc0001fffe0003ffff0007fffe0023f7ff1047c8ff80e39d7fc5c119238380951501451c300008a510000537b00009bdd0001dffb8003ffff0007ffff8003ffff0001ffff0000ff7f10017ffe20083e7470041c20e00e0001f00700";
 when "01000111101" => data <= 768x"ff80001fffc0011fffe0023fff70031ffff0023f5ff4071c8ffc2e1815745d143230082817400445a200004417000045b2022bfff77fffffffffffff775111f7ff0001ffff0001fffe0000ff7f10047ff820043ff060041fe0e0060201f00700";
 when "01000111110" => data <= 768x"ffe0001fffc0011fffe0031fff71011ffff0030e5ffc471c4ffc3e026530141426000222444000444400002244111177efbfffffffffffffffeeaefff7100177fe0000ffff00007ffe0000ff7c40047ff820003ff0400417c0e0020301c00701";
 when "01000111111" => data <= 768x"ff80018fffc10107ffe0018fff7101077ff8078e5f7c1f05c0200e035d0005118c8000318c00001188000031dc011131dfbffffffffffffffffeaafffd00007ffe00007ffc00007ffc00003f7c400077f840023fd040060780c0020301c00301";
 when "01001000000" => data <= 768x"ffe00083ffc001c7fff003837ff417c73ff83f80045016059800028811000114180000181000001c380000181101111dbbbffffffffffffffffeaefffd000077f800003ffc00001ff800003ff040011ff880021fc0c001078080030101c00100";
 when "01001000001" => data <= 768x"ffe000e1fff405c1fff80fe17f71174100e007005040004432000086310000043000000e700000047000000e7111111ffbbfffffffffffffffeeaebff100001ff800001ff000001ff000000ff100011fe080000fc10001050180018001000100";
 when "01001000010" => data <= 768x"fff803f0fff417f0fbe00f8011000101e0000001440000456000000240000007e0000003c0000007e000000770011117f3bffffffffffffffffeaeaf71000017e000000fc0000007e000000741000007e1000007410000050300008007000040";
 when "01001000011" => data <= 768x"fff007f8554001c4000000804400001580000002c000000180000001c000000180000003c0000001c000000340111107ebbfffffffffffffffeeeeafd100000780000003c0000001800000030000000182000003040000410600004004000040";
 when "01001000100" => data <= 768x"020000c040000051880000011000000100000000000000000000000000000001800000010000000180000001c00111118bbffffffffffffffffeaeab11000001000000000000000100000000000000000000000004000000080000001c000010";
 when "01001000101" => data <= 768x"2000000010000000000000000000000000000000000000000000000000000000000000000000000000000000011111112bfffffffffffffffeaa0808000000000000000000000000000000000000000000000000100000000000000010000010";
 when "01001000110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001155555bfffffffffdd555580000000000000000000000000000000000000000000000000000000000000000000000040000000";
 when "01001000111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000315555557ffffffff5555555500000001000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01001001000" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000085557577fffffffff5500001700000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01001001001" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000c057777f75fbaa2afe0000005f00000003000000010000000000000000000000000000000000000000000000000000000000000000";
 when "01001001010" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000000100000283577777d7a20003ff0000005f0000000f000000010000000300000001000000010000000000000000000000000000000000000000";
 when "01001001011" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000030000001f00aaae3f5757577f200003ff0000007f0000000f000000170000001f00000017000000070000000700000007000000070000180700001407";
 when "01001001100" => data <= 768x"0000000300000001000000010000000100000000000000000000000000000000000000380000007c00aab8fc555557fc000003fe0000017c0000007e0000007f0000003e0000001c0000003e0000001f0000203f0000541f00000c3f0000017f";
 when "01001001101" => data <= 768x"000000100000001000000008000000050000000300000001000000000000000000000020000001f00afefbf015555ff0000003f0000001f0000001f800000170000000f0000000f0000000f800004170000020f8000015f5000007ff00000375";
 when "01001001110" => data <= 768x"00000000000000400000002000000011000000110000001f000000000000000000000080000005c00affefc015555fc0000007c0000007c0000003c0000001c0000003c0000001c0000003e00000534700001bfe000007d000000fe0000177f0";
 when "01001001111" => data <= 768x"00000000000000070000000f0000001f0000000f000000570000000800000000000002000000070002ffff0015115f0000000f800000070000000f80000007000000070000010704000087980000777000001f8000015f400003ffe000017fd5";
 when "01001010000" => data <= 768x"0000000000000000000000380000007c0000007e0000007f0000003e0000000000000000c0045c0082fefe0045111f00c0000e00c0001f00c0000e00c0001f00c0000e00c0015f508000efc000001f0000003f0000057f400000ff28000177c0";
 when "01001010001" => data <= 768x"0000000000000140000001e0000001f0000001f80000015c0000002e000000010000000050155c0020eefc0071111c00f0001e0070001c0060001c0070001c0060021c0050015d4080007e0000017d000003ff800005ff400001ff000001f700";
 when "01001010010" => data <= 768x"00000f000000070000000f80000005c0000000e00000005c00000008000000000000000010055c0030eafc0011007c0038003c0070001c003000180010001c003002398050015d000000780000057d000007fe800001fc000003ff000007ff00";
 when "01001010011" => data <= 768x"00003e00000014000000020000000100000001e0000000500000000800000000000000001015500018eafc0011007c00180038001c001c00180038001c00310018023b00500174000000f8000005fd000001fc000001fc000003ff000005ff00";
 when "01001010100" => data <= 768x"0000f80000005c00000006000001070000000180000000500000000000000000000000001c05540008eaf8001c017c00180038001c007000080038001c00710018023a00540174000000f8000005f5000003fc000001fc000003fe000005fc00";
 when "01001010101" => data <= 768x"0003f0000001dc000001ce000001070000000380000000400000000000000000000000000c055400082afa001c117d001c0038001c0070000c0038001c00710018023a00500170000000f8000005f5000003f8000001fc000003fe0000057400";
 when "01001010110" => data <= 768x"0000f80000005c00000004000000070000000180000000400000000000000000000000001c55540008eafa001c007d001c0038001c0070000c0038001c00710018023a00500174000000f8000005f5000003fc000007fc000007fe000005fc00";
 when "01001010111" => data <= 768x"0000700000005c0000000400000003000000010000000040000000000000000000a000001c555000080078001c007400180038001c007000080030001c00710018023a00500174000000f8000005fd000003fc000001fc000007fe000005fc00";
 when "01001011000" => data <= 768x"000ff000000474000000240000010100000001000000000000800000015000000000e0001c01f0000800f0001c0074001800e0001c0040000800ec001c1170002803e0005001f4000007f8000015fc000003fe000007fc000007f80000041000";
 when "01001011001" => data <= 768x"00007000070074000f80780007c171000380000000400000000380000017c000000380001c01c0000803e0001c0350001803b0001c01c000080b80001c07d400280fe0005057f0000007f800000770000007e00000054000000c200000103000";
 when "01001011010" => data <= 768x"0000780000005c0000003e0000001c0000000000c0450000e00f800070170000200700001c070000080f80001c071000180f20001c4740000c0f80001c07d000281f8000505fc000001fe000001fd000000f8000000440000008400000004000";
 when "01001011011" => data <= 768x"0000238000001fc000000f80010005000000000000570000001f000000170000000e00001c1f0000080e80001c1440001c2e80001d5700000c0f0000141f5000286f8000505fc000001fc000001f4000000b0000000d00010008800000110000";
 when "01001011100" => data <= 768x"000023f004001ff002000ee00100000000020000005f0000001e0000001c0000001e00001c1d0000081c00001c1c40000c2e80001c5f00000c3f8000155f1000281f8000501fc000001f8000001f000000090000001900000008800000110000";
 when "01001011101" => data <= 768x"000023e004001ff000000af801000071001a0030001f0000001e0000001c0000001c00001c1c0010081c00001d1c40000c2f80000c5f00000dbea00015170000383f0000501f0000003f80000015000000090000001100040008800000110000";
 when "01001011110" => data <= 768x"00002000040017d0000008f801000071000f0070001f0050001e000000140000001e00000c1c0040081e00001d1440000c2f80000d7f00000c9f8000141f5000383f0000507f0000003f0000001d000000090000001100000008800000110010";
 when "01001011111" => data <= 768x"000020f0000017f0000000f000000050000080000007c0000007800000070000000300000c07c000080fc0001c1700000c1f00000c1750000cff8000145f5000083fa000507f0000007f8000001f000000088000000d80000008800000104010";
 when "01001100000" => data <= 768x"000020e0000015f0000000e00000014000000000000140000003c0000003c000000380000c05c4000c07e0001c0750000e2b90000c1d54000c7f82001417c1000807e0005017c040003fe020001fc110000f8000000c40050008800000104000";
 when "01001100001" => data <= 768x"00000000000055c0000009e0000001c000000080000540000007c0000007c000000380000407d0000c07e000140770000e2b30000c1f54000cff80001457d1000807f8005007f040000ff0200007c010000b8000000c40040008800000104001";
 when "01001100010" => data <= 768x"00000000000055c0000003e0000001c0000000800007c0000007800000070000000300000407c0000c0fc0001c0750000e2b30000c1f54000c3f80001457d100080ff0005007f040000fe00000174010000a8000000c40040008800000104000";
 when "01001100011" => data <= 768x"00000380000007c0000003e000000100000080000007c000000f800000070000000300000407c0000c0fc0001c0750000c2b30001c1f50000c2f80001d47d100080f8000500fc100000fe00000174010000a8000000c40140008800000104000";
 when "01001100100" => data <= 768x"00000f80000005c0000000e0000000000003800000070000000f800000071000000700000c07d000080f30001c1710001c0f20001c1f50000cef88001d07d400280f8800501fd500000fca000017150000088a00000c454000088a8000105550";
 when "01001100101" => data <= 768x"00030f0000150540000a80e000154000002be0000057d400000fa000005750010027f8000c5f4400080f00001d5701001c2f22001c5f40000caf80001d57d010280f8000505fc000000fc0000017000000088000000c40000008800000104000";
 when "01001100110" => data <= 768x"00003f0000007d54000038e0000111550003802200075555000f0eaa000755550007803a1c1f0015080f00021c5700011c1f80001c1f00000c2f80001d57d0002a0f8000501fc000000fc0000005000000088000000c40000008800000104000";
 when "01001100111" => data <= 768x"00003f0000001d40000000c0000001000002800000070400000f3e000007c400000788001c0f1400080f38001c5735001c1f20001c1f55000c2fc8001d57d5103b0fe000541fd540001fc0000015000000088000000840000008800000105000";
 when "01001101000" => data <= 768x"00000b0000000140000000c00000404000038000000785000007be0000075400000790001c075000080bc0001c570000180f00001c1f0000083f80001c57c0001b8f8000541fc000001fc000011f400000088000000c40000008800000104000";
 when "01001101001" => data <= 768x"00000780000005400000002000004010000380000007c50000038f80000175000003a80014071000180fe00010174000181b00001c1f0000181f80001c574000198fa000551fd000081fc000001f4000000f8000000c40000008c00000104000";
 when "01001101010" => data <= 768x"000001e0000001f0000000e0000040140001e0200001c5400003ef800001f5100003e6001007d400180fa00010574100183b80001c170000181f800018771000188fc000551fd000081fc800101f4100001fe000001fc0000008c00000184000";
 when "01001101011" => data <= 768x"0000003e0000001d0000001e000111050001e0080001c0500003e3e0000157400003fb001007c400180f880010475000382be0001c17c000180f80001017c000382f8000514fc0008e0fe800151f4400003fe000001ff000000fe00000154000";
 when "01001101100" => data <= 768x"0000000f0000000100002000000170010003e0010001c0050003e00c0001d1500003fbe01007d5c0180fc38010174500380bb8001c17d000180b80001017d000383fc000105fc000f38fe000171fd400381fe200001ff000001ff000041ff000";
 when "01001101101" => data <= 768x"00000000000010000000b000000170000003e0000007f0000003e0000001c0010003f8021007fdf0180feee011074140388bc6001c5fdc00183be0001017c000380fc000101fc000a8efe000515f74003e1ff600541ff100001ff8000017f000";
 when "01001101110" => data <= 768x"00000000000010000000d0000001f0000003e0000007f0000003e0000001c0010003f0031007fc44380ffff81107d570380bc3a01d5fc500382bd800101ff000380fe0001007c000283fe000517f7000238ffe001d1ff540781ff800101ff000";
 when "01001101111" => data <= 768x"00000000000010000001f000000370000003e0000007f0000003e0000001c0000003e0011007f005380ffe8811075770380bc0e01d1fc540388fce001057d000381fe0001007c000280fe000507f740000eff600171ff1403c1ff800501ffc00";
 when "01001110000" => data <= 768x"00000000000110000001f000000770000003e0000007d0000007e0000001c0000003e0001007f005180ff8081017dd51380bc3c01d1fc5c0388fce001057d400381fe0001007c000380fe000501f740000fff380155ff1400e1ff800701ff900";
 when "01001110001" => data <= 768x"00000000000110000003e000000770000007e0000007c0000007c000000140000003c0001007d004180fe00a101f7511380fbf801c1fc7003b8f8f001157d410383fe0001007c000380fe000511ff500007ff3a015dff0400e1ff800141ff800";
 when "01001110010" => data <= 768x"00002000000150000003e000000770000007e0000007c000000fc00000074000000780001007c004180fe00e111f7054380fbe801c1fc7003a0f8f0011575500383fe0001017c000380fe8005017f500003ff0a011dff0000f1ff800141ff000";
 when "01001110011" => data <= 768x"00002000000150000003e000000760000007e0000007c000000fc00000070000000780001007c000180fe00c111fc054381ff8801c1fd5043e0f8e0011575500183fe0001417c000380fe800501ff740003ff00011dff000039ff800151ff000";
 when "01001110100" => data <= 768x"0000207f0004417f000fe0ff001f417f003fc0bf001f415f003f803f0017105f001f003f001f4057003f800b003fc075003fe0b0005f5d10003f0e00141f1c0003bf3800017fc000003f8000013ff000003f8f00007fc10000ffc00001ff4000";
 when "01001110101" => data <= 768x"003ffffe001ffffd003ffff8001f7f75001ffffe001ffffd003fffff007fffff003fffff001fffff001fffff001f7f7f003fffff001ffffd000fffff0017f7f70002ff8300017d0700007e0700017f170000ff0f00017c170000fc0f00017417";
 when "01001110110" => data <= 768x"00fff82001fffc4001fffc8801ff751501fffb0a01fff51503fff88203fff90503fffa0f05fffc5707ffffce077f7fd00ffffff01ffffff40fffffe007f7f7d007fff3f005ffd7d0007e87e0000007c000000fe0000007c000000fe0000017f0";
 when "01001110111" => data <= 768x"001f8000001fc000007fe000007f514000ffe20001ffd44003ffe88007ff515107ffe22007ff445507ffe03e177ff5551ffff8e01fffd5403ffffae01ffff5701ffffa201fffd57007ff30300155107000003070000050700000382000007030";
 when "01001111000" => data <= 768x"0000000000050000000f8000011fc000003fc000005fd500007fe20001ffd54003fff80007ff554407ffe820077f51550fffe2301ffff5441ffff3001ffff5700ffff8f00fffd41007ff30380155301100003030000070100000301000007010";
 when "01001111001" => data <= 768x"00000000000000000000000001070000000fc000001fc000001fe0000077d50001ffe00001ffd54003ffe000037f515503ffe23807fff5540ffff08017fff5512ffffa6817ffd45c23ffb00c7155101c200030084000701c6000300870007004";
 when "01001111010" => data <= 768x"00000000000000000000000001074001000fe000001fc000000fe000005ff10000ffe20001ffd54003ffe800017f755503fff02807fff5540ffff88007fff5100ffffa321ffff4141bfff8021177100738003003100010071800380210003001";
 when "01001111011" => data <= 768x"0000000000000000000000000107c001000fe000000fc000000fe000007ff10000fff20001fff44003ffe800037ff55103fff80207fff5540ffff8a81ff7f1400ffffa000ffffd040ffff8001dff5001380010001c0010000800380018001000";
 when "01001111100" => data <= 768x"0000000000000000000280000007c000000fe000001ff000003fe000017ff10103ffe20007fff54007ffe880077f75110ffff8021ffff5541ffff8381ffffd503ffffe001ffffd011ffff8021f7ff0001fbf30001c0010003c0030001d003000";
 when "01001111101" => data <= 768x"0000000000140000003e0000007f4000007fc000017fc0000fffe00017f7c5003fffe8007fffd5007fffe2007f7f5511fffff220fffff454fffff820f7fff550fffffa00fffff400fffff8007f7fd0003fffc0001d55c0001c00c0007401c000";
 when "01001111110" => data <= 768x"1f8000005fd000003ff800007f7d0000fff80000fffc0400fffc0000f7fd5000fffa0000fffd4000fff880007f7d0000ffff0000ffff1500fffe0c00ffff7000ffffa000ffff0000fffe00007f7c0000fff800007d4000007ee0000075700000";
 when "01001111111" => data <= 768x"e0000000c0000000e000000050000000f8000000d5000000cf800000d7c00000ffe00000fff00000fff000007f700000fff00000fff00000ffe00000fff00000fff00000ffc000007fe000007f7000007fe000007ff00000fff000007ff00000";
 when "01010000000" => data <= 768x"00000000000000000000000007f0000007f8000007fc00000ffc000017fc00003ffe00001ffc00000ffe00001f7c00003ffc00007ffc00003ffc000017f400001ffc00001ffc00001ffc00001f7f00003ffe00007fff00073ffe000e77f7001c";
 when "01010000001" => data <= 768x"000000000000000003a0000007f000000ff800001ffc00000ffc00001ffc00003ffc00001ffc00000ffc00001f7c00001ffe00001fff00001ffe000017f400001ff800001ffc00003ffc00003f7c00003ffe00007fff00007ffe00007ff70000";
 when "01010000010" => data <= 768x"00000000054000000fe000001ff000001ff800001ffc00003ff800007ffc00007ff800001ffc00001ff800001f7c00003ffe00001ffd00000ffc00001ff000003ff800007ffc00003ffc00007f7c00007ffe00007ffc00007ffe00007ff70000";
 when "01010000011" => data <= 768x"0000000005c000001fe000001f7000003ff000007ff00000fff80000f7f000007ff800007ff000003ff800007f7100003ff800005ffc00001ff800007ff000007ff000007ff40000fff800007f7c0000fffc0000fffc0000fffe0000f7ff0000";
 when "01010000100" => data <= 768x"01000000150000003f8000007f4000003fe000007ff00000fff00000fff00000fff000007ff000007ff000007f700000fff00000fff000003ff800007ff00000fff000007ff00000fff800007f7c0000fffc0000fffc0000fffe0000f7ff0000";
 when "01010000101" => data <= 768x"01000000010000000f8000001fc000003fe000007ff000007ff000007ff00000fff000007ff000007ff000007f700000fff00000fff00000fff0000017f000007ff000007ff40000fff800007f7c0000fffc00007ffc0000fffe000077f70000";
 when "01010000110" => data <= 768x"0180000005c000000fe000001f7000003ff800001ff800003ff800007ff000117ff800005ff000003ff800007f7000007ff8000077f400000ff800001ff000003ff800007ffc00003ffc00007f7d00007ffe00007fff00007ffe000077ff0000";
 when "01010000111" => data <= 768x"0080000005c000000ff000001f7100001ff800001ffc00003ff800007ffc00003ffc00001ffc00001ffc00001f7c00003ffc00001ffc00000ffc000017fc00001ffe00001ffc00003ffe00001f7f00003fff00003fff00003fff000037ff0000";
 when "01010001000" => data <= 768x"0000000001c0000007e00000177000000ff800001ffc00000ffc00005ffc00003ffc00005ffc00000ffe00001f7400000ffe00001fff00000ffe000017fc00000ffe00001fff00000ffe00001f7f00001fff00001fff00000fff80001fff0000";
 when "01010001001" => data <= 768x"000000000040000000c0000007f0000007f8000007fc00000ffe000017fc00013ffe00001ffc00000ffe0000077f00000ffe00000fff00000fff000017f5000007fe000007ff00000fff0000077f00010fff00000fff40000fff800007ffd000";
 when "01010001010" => data <= 768x"000000000040000400e00000077c000007fe000007fc00000ffe000017ff00003ffe00001fff000007fe0000077f000007ff000007ff00000fff000007ff100003ff000007ff000007ff8000077f000107ff800007ffc00007ff800007ffc000";
 when "01010001011" => data <= 768x"002000000070000001fc00000377000003ff000007ff000007ff000017ff00001fff000007ff000003ff000007ff000007ff000007ff000003fe000001ff000003ff800007ff000007ff8000077fc00007ff800007ffc00007ffc00007ffc000";
 when "01010001100" => data <= 768x"00300000017c000001fe0000017f000003ff800005ff000003ff800017ff000007ff800005ff000003ff8000077f400003ff800007ffc00003ff800001ff000003ff800005ffc00003ffc00007ff400003ffe00007ffc00007ffe00017ff4000";
 when "01010001101" => data <= 768x"00080000001c0000007e0000017f000101ff800001ffc00001ff800005ffc00007ffc00005ffc00001ffc000017fd00003ffc00007ffc00003ffe000017f400001ff800001ffc00003ffc000037f400003ffe00007ffc00007ffe00007ffc000";
 when "01010001110" => data <= 768x"00080000001c000000fc0000017f000103ff000001ff000003ff800003ff000007ff800005ffc00003ff800001ffc00003ffc00001ffc00003fee00001ff100003ff800001ffc00003ff8000077fc00007ffc00007ffc0000fffc00017f7c000";
 when "01010001111" => data <= 768x"00080000005c000001fc0000037f000003ff000007ff000007ff00001fff00000fff000007ff000003ff000007ff000007ff800007fdc00003fc000007ff000007ff000007ff00000fff8000077f00000fff800007ffc0000fff80001fffc000";
 when "01010010000" => data <= 768x"000000000150000003f80000477c000007fe000007ff00000ffe00001fff00000fff000007fd00000ffe0000177f00000fff000007ff000007fe000017fe00000ffe00001fff00000fff00001f7f00001fff00001fff00001fff80001ff70000";
 when "01010010001" => data <= 768x"000000000010000001f8000007fc000007fe000017fc00000ffe000017fe00001ffe00000fff00000ffe00001f7c00001ffe00001ffc00000ffe000017fd00000ffe20001ffc40001ffe60001f7f40003ffe60001fff40003fffc00037f74000";
 when "01010010010" => data <= 768x"000000000010000000b0000007f000000ff800000ffc00000ffc000017fc00003ffe00001ffc00000ffe00001f7c00001ffc00001ffc00003ffc000017fc00101ff820001ffc70003ffe60001f7f70003ffe60007fff40003ffe60007ff74000";
 when "01010010011" => data <= 768x"000000000040000003e0000017f000001ff800001ffc00001ffc00007ffc00003ff800005ffc00001ffc00001f7d00003ffc00001ffc00003ffc000017f000103ff8f0001ffcf8003ffcf8007f7c71003ffef0007ffc70007ffee0007ff77000";
 when "01010010100" => data <= 768x"00000000054000000fe000001f7000003ff800001ff000003ff800007ff00000fff800005ffc00003ff800007f7000003ff800007ffc00003fec000057f150007ff3f8007ff7fc007ffffe007f7ffc00fffff8007ffdfc00fffff8007ff7f000";
 when "01010010101" => data <= 768x"00000000058000003fc000003ff000003ff000007ff00000fff00000fff10000fff000007ff400007ff000007f7100007ff800007ff000003ff8000077f15000fff3f8007fffff00ffffff807f7f7fc0ffffff80ffffff00fffffe00fffffc00";
 when "01010010110" => data <= 768x"00000000010000000b8000001f4000003fe000007ff000007ff000007ff04000fff000007ff040007ff000007f700000fff00000fff00000fff0000057f150003fe3f8007ff7ff00ffffff807f7f7fc0ffffffe0fffffff0ffffffe07f77f750";
 when "01010010111" => data <= 768x"00000000010000000f8000001ff000003ff000001ff000003ff800007ff04000fff020007ff010003ff000007f700100fff80000fff000006ff8000017f000003ff820007ffdfc007fffff007f7f7fc07fffffe07ffffff0ffffffe077ffffd0";
 when "01010011000" => data <= 768x"0080000005c000000fe000001f7000001ff800001ffc00003ff800007ffc00007ff800001ffc00001ff800001f7c00003ffc000077fc00000bf8000017fc00003ffc00001ffc00003ffe00007fff50003ffffe007fffffc03fffffe077fffff0";
 when "01010011001" => data <= 768x"0080000001c0000007e00000177000000ff800001ffc00001ffc00007ffc00003ffc00001ffc00000ffc00001f7c00101ffe00001ffe00000ffe000017fc00001ffe00001ffc00001ffe00001f7f00001fff00001fff00001fffa80017f7ff00";
 when "01010011010" => data <= 768x"000000000040000000c0000007f100000ff8000007fc00000ffc000017fc00003ffe00001ffc04000ffe0000077d00050ffe00000fff00000fff000017f4000007fe000007ff00000fff000017ff74000fffff001fffff400fffffc017ffff70";
 when "01010011011" => data <= 768x"000000000040000000e0000001f0000007fc000007fc00000ffe000007f500001ffe00001ffe04000ffe0000077f000007ff000007ff00000fff800017fd000003fe000007ff500007fffe0007ff7f000fffff8007ffffc00fffffe007fff7f0";
 when "01010011100" => data <= 768x"000000000040000000f8000007fc000003fe000007ff000007fe000017ff00001fff000017ff000007fe0000077f000007ff000007ff00000fff000003ff000003ff000007ff500007fffe0007ff7f0007ffff8007ffffc007ffffe007fff7f0";
 when "01010011101" => data <= 768x"002000000074000001fe0000017f000003ff000007ff000003ff800017ff00000fff800007ff000003ff8000077f000007ff800007ff000003ff800001f7000003ff800001ffc00003ffc000077fd40003ffff0007ffffc007ffffe007fffff0";
 when "01010011110" => data <= 768x"00080000005c000000fe000001f7000003ff800001ffc00003ff800007ffc00007ff800005ffc40003ff8000017fc00003ffc00007ffc00003ff80000177000001ff800001ffc00003ffc000077fc00003ffe00007ffdd0007ffffc007fffff0";
 when "01010011111" => data <= 768x"0000000000040000000c0000017f000001ff000001ff000003ff800001ff000003ff800007ffc00003ff8000017fc00003ffc00001ffc00003ffe00005f5400001ff800001ffd40003fffe00077f7f4003ffffc007ffffc007ffffe007fffff0";
 when "01010100000" => data <= 768x"00000000001c000000fc000003fc000003fe000007ff000007ff000007ff000007ff800007ff000007ff0000077f010003ff800007fd400003f800000375000003ff000007fffc0007ffff00077f7f400fffffe007ffffd00ffffff017f5f7f0";
 when "01010100001" => data <= 768x"001000000150000003f80000077c00000ffc00001ffc00000ffe00001ff700001ffe00001ffc04000ffe0000077f00000fff000007f400000ff8000007fc000007fe000007ff54000ffffe001f7fff000fffffc01fffffc00ffffff01ff7f7f0";
 when "01010100010" => data <= 768x"002000000050000002f0000007f100000ff800001ffc00001ffc00001ff500001ffe00001ffc00001ffc00001f7c04001ffc00001ff400001fe0000017f400000ffe00000ffc00000ffe00001f7f00011fff00001fff55001fffff801ff7fff0";
 when "01010100011" => data <= 768x"000000000040000000600000057000000ff000001ff800001ff8000017fc00001ffe00001ffc00001ffc00001f7c04001ff800001ffc00003fe8000077f000008ffc20001ffdfc001fffff801f7f7fc03fffffe05ffffff03ffffff07ff7f7f0";
 when "01010100100" => data <= 768x"000000000040000000c00000177000001ff000001ff000003ff800003ff400003ffc00001ffc00003ff800001ff001001ff802001ff400003fe000001ff000007ff820005ffdfc003fffff007f77ff003fffffc07fffffc07fffffe07ff7f7f0";
 when "01010100101" => data <= 768x"00000000004000000fc000001f7000003ff000007ff000007ff800007ffc00003ff800007ff000003ff800003ff001003ff000001fd000003f80000037f000003ff800007ffdf4007ffffe007f7f7f007fffff807fffffc0ffffffe07ff7f7f0";
 when "01010100110" => data <= 768x"00000000010000000f8000007fc000007fe000007ff00000fff800007ff400007ff000007ff000007fe002007f4001007fe000007fc000007f8000007ff00000fff000007ff00000fff800007f7c0000fffff800fffffd00ffffff80ffffffc0";
 when "01010100111" => data <= 768x"0000000000000000008000001fc000007fc000007fc00000ffe00000fff00000fff000007ff00000ffe002007fc00100ffc000007fc00000ff80000077500000ffe000007ff00000fffaa0007f7ff400ffffff00ffffff00ffffffc0ff77f740";
 when "01010101000" => data <= 768x"00000000004000000080000017c000003fe000007fc00000ffe000007ff400007ff800007ff000007fe002007f4001007fe000007fc00000ff800000575000003ff000007ff150007ffffc007f7f7f007fffff807fffffc0ffffffc07ffff7c0";
 when "01010101001" => data <= 768x"000000000050000003e000001ff000003ff000007ff000003ffc00007ffc00003ff800001ffc00003ff002001ff000003ff000007fc000007fe0000057f00000bff800001ffdd0003ffffe003f7f7f003fffff807fffffc03fffffc077fff7c0";
 when "01010101010" => data <= 768x"000000000044000003e0000017f000001ff800001ff000003ffe00001ffd00003ffc00001ffc04001ff800001f7000000ff000001fd000001fe00000177c00003ff800005ffc00001ffe00001f7f74001fffff001dffffc03fffffc01dfff7f0";
 when "01010101011" => data <= 768x"000000000000000000200000057000000ff800001fdc00001ff800001fff00001ffe00001ffc04000ff800001ff100000ff8000007f000000fe00000177400000ffc00001ffc00000ffe00001f7f00000fffba001fffff400fffffc01ffff770";
 when "01010101100" => data <= 768x"0000000000000000002000000170000003f8000007fc00000ffc00001ff700001fff00001ffe00000ffe0000077c00000ff8000007fc00000ff80000077400000ffe200007fdfc000fffff00077f7f400fffffe007ffffe00fffffe007fffff0";
 when "01010101101" => data <= 768x"0000000000100000003000000170000007f8000007fc00000ffe00001fff00000fff000007ff040007fe0000077c000007fe000007fc000007f8000007f500000ffe20001ffffd000fffff80077f7fc007ffffe007fffff007fffff007fffff0";
 when "01010101110" => data <= 768x"000000000010000000f80000017c000007fe000007fd00000fff800007ff00000fff000007ff000007fe0000077f000003fe000007f4000007f8000007f7000007ff000007ff54000fffff80077f7fc007ffffe007fffff007fffff807fffff0";
 when "01010101111" => data <= 768x"000000000050000000fc000001fc000003fe000007ff40000fff800007f7100007ff800007ff000003fe0000177f000003fe000007fc000003fe000007ff000003ff800007ffc00007ffc000077f400003ffe00007ffdfc007fffff807fff7fc";
 when "01010110000" => data <= 768x"000000000000000000080000007c000001fe000005ff000003ffc00007ff400007ff800007ffd00003ff8000017f000003ff000001ff000001fe000001f5000003ffb80001ffff0003ffffc0077f7f7003fffff007fffff007fffff807fff7f0";
 when "01010110001" => data <= 768x"0000000000100000003000000174000003fc000007fc00000fff800017ff00000fff000007ff100007fe0000077f000003fe000001fc000003f8000001f5000003ffba0007ffff4007ffffc0077f7f700ffffff007fffff00ffffff817ffffd0";
 when "01010110010" => data <= 768x"000000000040000001f0000007f100000ff800001ffd00001fff000017f700001ffe00000ffc00000ffc0000077c000007fc000007f0000007f8000017fd00000ffe380007ffff000fffffc01f7f7f500ffffff01ffffff00ffffff81ffdf7f0";
 when "01010110011" => data <= 768x"000000000040000000e0000007f100000ff800001ffc00001fff00001ff500001ffe00001ffc00000ff800001f7d00000ff800000fd000000fe000001ff500000ffe00001fff00001ffe00001f7f55001fffff801ffffff01ffffff81ffff7f0";
 when "01010110100" => data <= 768x"000000000040000000200000057000000ff000001ff000001ff8000017ff00003ffe00001ffc00000ff800001f7000001ff800001ff000001fe00000177000003ffe00005ffd54003ffffe001f7f7f403fffffe01ffffff03ffffff037f7f7f0";
 when "01010110101" => data <= 768x"000000000040000000400000077000000ff000001ff000003ff8000077fc00003ffc00001ffc10001ff800001f7000001ff000001ff000001fe000001fd000003ff8b0007ffdfc003fffff003f7f7f403fffffc07fffffc07fffffe07ff7f740";
 when "01010110110" => data <= 768x"00000000000000000280000017c000003fe000007ff00000fff800007ffc00007ff800007ff010003ff000007f7000003fe000001fc000003f800000375100003ff8a0007ffffc007ffffe007f7f7f007fffff807fffffc0ffffffe07ffff7f0";
 when "01010110111" => data <= 768x"00000000010000003f8000007f400000ff800000ffc00000ffe80000ff701000fff01000fff01000ffe00000ffc00000ffc000007fc00000ff80000077500000ffe00000fff00000fff800007f7f7400ffffff00ffffffc0ffffffc0fffff7f0";
 when "01010111000" => data <= 768x"0000000004000000fe000000ff000000ff000000ff000000ffa00000fff00000ffe02000ffc00000ffc000007f000000ff800000ff000000ff000000fd000000ff800000ffc00000ffe000007f700000fff00000fffd5400fffffe00ffffff40";
 when "01010111001" => data <= 768x"00000000040000002c00000074000000fe000000ff000000ff000000ff500000ffe04000ffc04000ffc000007f000000ff000000ff000000ff000000f7000000fe000000ff400000ffc3e0007f577d00ffffff00ffffff40ffffffc0fff7f7c0";
 when "01010111010" => data <= 768x"0000000050000000fc000000ff000000fe000000ff000000ff800000f7f00000ffe08000ffc44000ff8000007f010000ff800000ff000000ff000000ff000000fa000000ffc00000ffc00000ff455000fffffe00ffffff00ffffff80fff7f7c0";
 when "01010111011" => data <= 768x"2000000070000000f8000000fc000000fe000000ff000000ffe00000ffc10000ff800000ffc00000ff8000007f010000ff000000ff000000ff000000ff000000f8000000fd400000ffc000007f400000ffe00000ffd00000fff00000fffff400";
 when "01010111100" => data <= 768x"80000000c0000000e000000070000000f8000000fc000000fe800000ffc10000ff800000ff000000ff8000007f000000ff000000ff000000ff000000ff000000fe000000fc000000f80000007f400000ff800000ffc00000ffc00000ffd00000";
 when "01010111101" => data <= 768x"00000000000000000000000040000000e0000000f0000000f8000000fd000000ff800000ff000000ff0000007f000000ff000000fd000000fe000000ff000000fe000000fd000000fe0000007c000000f0000000f5000000ff800000f7c00000";
 when "01010111110" => data <= 768x"0000000000000000000000000000000080000000c0000000e0000000f1000000ff000000ff000000fe00000077000000fe000000fc000000fc000000fc000010fc000000fc000000fc0000007c000000f8000000d0000000e8000000ff000000";
 when "01010111111" => data <= 768x"0000000000000000000000000000000080000000c0000000c0000000f7000000fe000000fc010000fe0000007c000000fc000000fc000000f8000000f0000010f8000000fc000000f800000074000000f0000000f0000000c000000040000000";
 when "01011000000" => data <= 768x"0000000000000000000000000000000000000000000000008800000074000000fc000000fc000000fc0000007c010000fc000000fc000000f8000000f0000000f0000000f0000000f000000070000000f0000000f0000000e0000000c0000000";
 when "01011000001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000008020000dc030000f8030000f0010000f8000000dc000000f8000000f0000000f0000000f0000000e000000071000000e0000000c0000000e0000000f0000000";
 when "01011000010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000400000002000000010000800100000000000000000000000000008000000000000000800000000000000000000000000000000000000000000000";
 when "01011000011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000400000002000000030000000300000001000000008000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01011000100" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000040000000f0000001700000007c0000007c0000000e000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01011000101" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000040000000f8000001fd000001ff000001fd00000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01011000110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000040000003f00000177000001fe000001fc000000f0000000400000000000000000000000000000000000000000000000000000000000000000000";
 when "01011000111" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000030000001f0000003e0000007c0000007c0000007c000000f8000001710000002000000000000000000000000000000000000000000000000000000000000";
 when "01011001000" => data <= 768x"000000000000000000000000000000000000000000000000000000000001c0000001e0000001c0000003c0000003c0000003c0000007c0000007c0000007c0000007800000050000000000000000000000000000000000000000000000000000";
 when "01011001001" => data <= 768x"0000000000000000000000000000000000000000000100000003000000071000000380000007c0000003c0000007c0000003e0000001c0000003e0000001c0000001e0000001c000000080000000000000000000000000000000000000000000";
 when "01011001010" => data <= 768x"000000000000000000000000000000000000000000040000000e000000070000000f0000000740000007c0000007c0000003e0000001f0000001f0000001f0000000f80000007000000020000000000000000000000000000000000000000000";
 when "01011001011" => data <= 768x"00000000000000000000000000000000000000000000000000000000001c0000001e0000001f0000000fc000000770000007f0000001fc000001fc0000007c0000003c0000001400000000000000000000000000000000000000000000000000";
 when "01011001100" => data <= 768x"0000000000000000000000000000000000000000000000000000000000500000007e0000007f4000003fe000001f7000000ffc000005ff000000fe0000007f000000020000000000000000000000000000000000000000000000000000000000";
 when "01011001101" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000028000000fd400000ffe000007ffd00003fff000007ff000000ff00000015000000000000000000000000000000000000000000000000000000000000000000";
 when "01011001110" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000001000000055400001fffe0001ffff0000ffff00005fff000002f800000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01011001111" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000002000000145400003ffe00017f7f0001ffff00007ffc00003f8000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01011010000" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000002000000545c00001bff00001fff0001fffe0001fff40000ff8000005500000000000000000000000000000000000000000000000000000000000000000000";
 when "01011010001" => data <= 768x"00000000000000000000000000000000000000000000000000000000001000000002080000145d00001bfe000017fc00003ff800017ff00000ffc000007d00000030000000000000000000000000000000000000000000000000000000000000";
 when "01011010010" => data <= 768x"000000000000000000000000000000000000000000000000000000000001000000020000001d7c00000bfc00001ffc00001ff800005ff000007fc000007f0000003e000000140000000000000000000000000000000000000000000000000000";
 when "01011010011" => data <= 768x"00000000000000000000000000000000000000000000000000000000000100000002000000057c00000ff80000177100000ff000001ff000003fc000001f4000001f0000001c0000000000000000000000000000000000000000000000000000";
 when "01011010100" => data <= 768x"000000000000000000000000000000000000000000000000000000000001000000030000000550000003f00000077000000ff000001ff000000fe0000017c000000f800000070000000200000000000000000000000000000000000000000000";
 when "01011010101" => data <= 768x"000000000000000000000000000000000000000000000000000000000001000000018000000140000003e00000077000000ff000000ff000000ff0000007f0000003e0000005c000000080000000000000000000000000000000000000000000";
 when "01011010110" => data <= 768x"00000000000000000000000000000000000000000000000000000000000040000000c0000000c0000002c000001f4000001fe000001ff000000ff800000770000003f0000001f000000000000000000000000000000000000000000000000000";
 when "01011010111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000600000006000000040000000600000177000003ff000001ff400000ffc000007fc000003f80000015000000000000000000000000000000000000000000000000000";
 when "01011011000" => data <= 768x"000000000000000000000000000000000000000000000000000020000000700000002000000070000000300000147100007ff200007ff700003ffe000017fc000003fc0000015400000000000000000000000000000000000000000000000000";
 when "01011011001" => data <= 768x"00000000000000000000000000000000000000000000000000002000000070000000300000005000000030000000710000ba798000ffff00007fff00001ff7000007fe0000055400000000000000000000000000000000000000000000000000";
 when "01011011010" => data <= 768x"00000000000000000000000000000000000000000000000000003000000050000000300000005000000038000000704000203a8001fd5f0000ffff800057ff00000ffe0000055400000000000000000000000000000000000000000000000000";
 when "01011011011" => data <= 768x"00000000000000000000000000000000000000000000500000003000000050000000100000005000000038000000704000207bc007fd5fc003ffff8001777f00003ffe0000055400000000000001000000000000000000000000000000000000";
 when "01011011100" => data <= 768x"00000000000000000000000000000000000000000000500000003000000010000000180000001000000038200000784002007be007f55fc007ffff80017f7f00003fff00001d5400000000000000000000000000000000000000000000000000";
 when "01011011101" => data <= 768x"0000000000000000000000000000000000000000000050000000b000000110000000100000001000000038000000713002003be01ff55fc00fffff800577ff0000ffff00005d7f00000000000000000000000000000000000000000000000000";
 when "01011011110" => data <= 768x"000000000000000000000000000010000000b000000050000000980000011000000030000001100000007818000071502a003be07ff55fc03fffffc01777f7c003ffff8001757f0000000e000000000000000000000000000000000000000000";
 when "01011011111" => data <= 768x"00000000000000000000000000017000000130000001140000001800000110000000380000017c040000f80800017170fa003bf0ffd55ff0ffffffe05ff7f7c00fffff8005d5ff0000003e000000140000000000000000000000000000000000";
 when "01011100000" => data <= 768x"0000200000017000000370000001150000023a000001100000023800000130010002780300007c070000f83e00017d7cfa003ff8ffd5fff0fffffff077fff7f07fffffe05d55ffc00000ff000000150000000000000000000000000000000000";
 when "01011100001" => data <= 768x"000670000004554000043800000410000004380000045c000004780000057c000000fc000001fc170000f8ff000037f7fa03fffefffffffcfffffff87ff7fff0ffffffe0f5dfffc08007ff8001017f0000001e00000004000000000000000000";
 when "01011100010" => data <= 768x"00103800001070000010380000107100001878000011fc000001fc000011fc010003f80f00057d7f00003fff00157fffbbfffffffffffffffffffffe7ff7fffcfffffff8fffffff0007fffe00017ffc00003ff0000005c000000000000000000";
 when "01011100011" => data <= 768x"00c07000004070000060f8000041f0000043f8000047f8000007f8000007f017000af0ff000077ff000bffff577ffffffffffffffffffffffffffffef7fff7f4fffffff8fffffff08fffffe005ff7fc000ffff800015f5000000000000000000";
 when "01011100100" => data <= 768x"0181f0000187f000018ff800011f7001001ff000005ff000003fe0030015f0570000e3ff00057fff2fffffffffff7f7ffffffffffffffffffffffffefffff7fcfffffff8fffffff0ffffffe07f7f7f003ffffe0005ff54000000000000000000";
 when "01011100101" => data <= 768x"0303f0000117f000021ff8000117f001013ff000017ff000003fe003001571570000e3ff0015dfffafffffffffff7f7ffffffffffffffffffffffffefff7f7fcfffffff8ffffffd0ffffff807f7f7f01fffff8005fff50000fa8000001000000";
 when "01011100110" => data <= 768x"0303f0000107f000020ff800011ff000023ff800015ff00000fff0000017f0170000e0ff0000d5ff000bffff577ffffffffffffffffffffffffffffefffffff4fffffff8fffffff0ffffff807f7f7d00fffff000ffff4000fffc000055500000";
 when "01011100111" => data <= 768x"0301f0000105f0000307f800031f7000023ff800015ff00000ffe000007ff0150003e03f0001d5ff0000efff0115ff7fbffffffffffffffffffffffffffffff7fffffffefffffffcfffffff07f7f7f50fffff000ffff4000fffe0000ff700000";
 when "01011101000" => data <= 768x"0601e0000701f0000203f80003077000020ff800041ff000023ff8000177f000003ff0030015f05f0000e3ff0001d7ff002fffff5d7ffffffffffffffff7fff7fffffffffffffffdfffffffc7f7f7f70ffffffe0ffffdd40ffff8000fffd0000";
 when "01011101001" => data <= 768x"0e03e0000401f0000600e0000701f0000203f8000407f800060ff800041ffc00020ff800015ff005003ff83f0001f17f0000ffff0555ffffbfffffffffffffffffffffffffffffffffffffff7f7f7f77fffffffefffffffcffffffe0ffffff40";
 when "01011101010" => data <= 768x"0c03e0001c01c0000c03e0001401f0000601f0000401f0000603f8000407f0000407f800041ffc00020ff80001177017003ff8ff0005dfff0001ffff15777fffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffefffffffc";
 when "01011101011" => data <= 768x"1801fe031c01f4001803e0001d03c0001c01e0001c01f0000c01f000040370000c03f0000407f0000c0ff800051f7001020ff003001ff05f003fe3ff0015f7f7002bffff55ffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffff";
 when "01011101100" => data <= 768x"3803e3a01c01e55d3803fe031003f0003803e0001c05c0001801e0001c01f0000c03f0000c07f000080ff000151f7001083ff000045ff000043ff003003fd05f003fe3ff0055dfff002fffff57ff7f7fffffffffffffffffffffffffffffffff";
 when "01011101101" => data <= 768x"3807c0001c05d4003801e380300175553803fe031005f4003803e0003001c0003801e0001c01f0001807f0001c1f7000083ff000187ff00008fff800107f700008fff00304fff05f00ffe3ff015f77ff003fffff5ffffffffffffffff7f7ffff";
 when "01011101110" => data <= 768x"3f87e0001c57c000380fc000700755003003e3807001c5d53003ff0f7003f4013003e0007005c0003801e0001001f0003803f0001c1ff000183ff8001077f00010fff80011fffc0008fff803057f701703fff3ff01ffffff00ffffff57ffffff";
 when "01011101111" => data <= 768x"3803e0001d07f00038cfe00071174001380780007005d4007003ef80700171d57003f38f7007fd017003e000700140003001e0007001f0003803f0001007f000381ff800107ffc0030fff80011ff7c0011fff80315fffc1703fff8ff07fff7f7";
 when "01011110000" => data <= 768x"000000005001c0003c03e0007d07700038a7e0007017c0007007c0007005f5007003e3807001f1d4e003ff8f70077f016003e0007001c0007001e0007001f0003003f0001007f400380ff800101f7000303ff800117ffc0010fffc0011fffc17";
 when "01011110001" => data <= 768x"00000000000000002003c0007407f0003e07f0007d47f000782fe0007017c000f003e0007001f500e003e1e0700171d5e003ff834007fc00e003e0007001f0007001f0007001f0003003f80031077400300ff800101ffc00207ff800117ffc00";
 when "01011110010" => data <= 768x"0000000000000000000000005001d0003803e0007d07f0007887e0007017c0007007c0007005d000e001ee00700171d0e003f1fe4007f705e003fe007001f0006000e0007001f0003003f00030077000300ff800301ffc00203ff800307ffc00";
 when "01011110011" => data <= 768x"000000000000000000000000110140003003e0007c07f0007a87f0007057f000700fe0007005c000e001f80070017540e003f0f86005f5c5e003ff007001f4006000e0007001f0007003f00070077000300ff800101ffc00203ff8003077fc00";
 when "01011110100" => data <= 768x"000000000000000000000000000100002003e0007c07f0007e07f0007157f000703fe0007007c000e001e0007001f500e003f1e06001f1d5e003ff837003f500e001f0007001f0007001f000700370003007f800101ffc00303ff8003077fc00";
 when "01011110101" => data <= 768x"000000000000000000000000000100002001a0007401f0003e03f0007147f0007823e0007017c000f003e0007001f501e001f3a07001f0d5e003fb837003ff01e003f0007001f0007000f0007001f0003003f8001007fc00380ffc00301ffc00";
 when "01011110110" => data <= 768x"000000000000000000000000000000000000a0007001f0003c03f0007507f0007823e0007017c000f003e0007001f501e001f3a07001f054e003fbc370037f016003f8007001f0007000f0007001f0003003f8001007fc00380ffc00101ffc00";
 when "01011110111" => data <= 768x"00000000000000000000000000000000000180005001f0003c03f0007507f0007823e0007017c000f003e0007001f500f001f3a07001f054e003fbc370037f016003fa007001f0007000f0007001f0003803f8001007fc003807fc001017fc00";
 when "01011111000" => data <= 768x"000000000000000000000000000000000001a0005007f0003c07f00075077000782fe0007017c000f003e0007001f500f001f3e07001f055e003fbc370037f006003f8007001f0007000f0007001f1003803f8001007fc001807fc001017fc00";
 when "01011111001" => data <= 768x"000000000000000000000000000000000003a0005007d0003807e0007507f000782fe0007017c000f003e00070017500f001f2e07001f055e003fbc07003f7006001f0007000f0007000f8007001f1003803f8001c07fc001807fc001017fc00";
 when "01011111010" => data <= 768x"000000000000000000000000000000000003e0005007e0007807e0007507c000782fe0007017c000f003f0007001f550f001f0fa7001f1c5e003ff807003f5007001f0007000f0007000f8007001f1003803fc001c07fc00180ffc001017fc00";
 when "01011111011" => data <= 768x"000000000000000000000000000140000003e0005007c0003c0fe0007557c000783fc0007007d000f003f8007001f5747003f8eb7001f5c1e003ff00700174007000f0007000f0003000f8003001f4003803fc001c07fc00180ffc00101ffc00";
 when "01011111100" => data <= 768x"000000000000000000000000000140000007e0005407c0003e0fe000715fc000703fc0007007f0007003fec07001f1757003f8c37003ff406003fe007001f0007000f0007001f0003001f80030017c003803fc001c07fc00080ffc00181ffc00";
 when "01011111101" => data <= 768x"000000000000000000000000000540000007e0007407c0003e0fe000715fc000782fe0007007f4007003fae07001f1757003fbc07003ff407003fc00700170007000f0007001f0003801f80010037c001807fc001c17fc00081ffc001837fc00";
 when "01011111110" => data <= 768x"000000000000000000000000000540000007e000740fc0003e0fe000715fc000780fe0007007f4007003fae07001f0777003fbc070037f007003f800700170003000f0007001f0003801f8001c077c00180ffc001c1ffc00083ffc001c77fc00";
 when "01011111111" => data <= 768x"00000000000000000000000000054000000fe000741fc0003e1fe000717fc000780fe0007007f4007003fae07001f0777003fbc070017f007003fc00700170003000f0007001f0003801f8001c077c00180ffc001c1ffc000c7ffc001c7ff400";
 when "01100000000" => data <= 768x"000000000000000000000000000140000007e000141fc0003e1fe0007d5fc000380fe0007007f4007802fae07001f0777001f8e070017f407001fe00700170003000780030007c003801fc001c077c001c1ffe001c5ffc000cfffc00157ffc00";
 when "01100000001" => data <= 768x"000000000000000000000000000170000003f0001c07f0003e8ff0001d57f0003803f0007c05fc003803fea070017c753800fe307801ffd03801ff8030007d0038003c001c007c001c00fe001c05ff000e0fff00045fff000e7fff00047fff00";
 when "01100000010" => data <= 768x"000000000000000000000000000074000001f8001d01fc000f83f8001f5774001e03f8001c01ff003c00ffe81c007f173c003f0e1c005f5c1c00ffe01c0077401c003e001c001f000e003f00150177000e03ff800707ffc0071fffc00777ffc0";
 when "01100000011" => data <= 768x"00000000000000000000080000001f0000003f0007007f000fe0fe001715ff000f01fe001f007fc00e003ff81f001fd51e001fe11e0017c70e003ffe1e0017d40e000f800f0007c00e000fc007001fc007003fe007007ff00380fff001c5f7f0";
 when "01100000100" => data <= 768x"000000000000000000000380000007c002001fe007c01fc007e83fc007c577c007803fc0074017f00f800ffe070007750f0007f8070007fc0f000fff070005f7078003f2070001f0078001f8070001fc038003f801c007fc01c00ffe01c01ff5";
 when "01100000101" => data <= 768x"0000000000000050000000f80100077c03a007f801f407fc03ef9ff801f15df003e00bfa07c001ff03c003ff07c0017f03c000ff07c001ff03c003bf07c0017f03c001ff01c0007f03c0003e01c0007701e000ff01e001ff00e003ff007017ff";
 when "01100000110" => data <= 768x"000000020000001f0000007f0150017f00f801ff01fd45ff00f8fbff01f0177f01f000ff01f0007f01e000ff01f0005f01e0003f01f0007f01e0006f01f0007701e0003f01f0001f00e0000f01f1001700f0000f0070001f0078003f0074017f";
 when "01100000111" => data <= 768x"00000003000000070060000f007d011f007f803f007c557f00fc03ff007c017f00f8003f00fc001f00f8001f01f1001700f8000701f0000700f8000d01f0001d00f8000f0070000700f800030078000100780001007c0005003c000700140017";
 when "01100001000" => data <= 768x"0000000000740007003f8007003fd007003f3f0f007f05df007e002f00770005007e0003007c000100fc0003007c0001007c0001007c000100fc0003007c0007007c0003007c0001007c0000007c0000003e0000001c0000003e0000001f0000";
 when "01100001001" => data <= 768x"003f8000001fd001003ffe00001fc575003f803f007f0005003f0000007f0001007f0000007f0000007e0000007f0000007e0000007f0000007e0000007f0000003e0000007f0000003e0000007f0000003f0000001f0000001f0000001f0000";
 when "01100001010" => data <= 768x"001ffffa001ff15f003fe003001f4000003fc000007fc000003f8000007fc000003f8000007fc000007f800000770000003f8000007f0000007f800000770000003f8000007f0000003f8000003f0000003f8000001fc000001f8000001fc000";
 when "01100001011" => data <= 768x"001ff800001ff800003ff800001ff000003ff000001ff000003fe000007ff000003fe000007fe000003fe000007f6000003fe000007fc000003fe0000077e000003fe000003fc000003fe000001fe000003fe000001ff000001fe000001ff000";
 when "01100001100" => data <= 768x"001fff00001fff00003ffe00001fff00003ffe00001ffc00003ffe000037f400003ffc00001ffc00003ffc00003ffc00003ffc00001ffc00003ffc00001ff400003ffc00001ffc00003ffc00001f7c00001ffc00001ffc00001ffc00001ffc00";
 when "01100001101" => data <= 768x"000ffff0001ffff0000fffe0001f7ff0001fffe0001fffc0001fffe0001fffc0001fffe0001fffc0001fffc0001f7fc0001fffc0001fffc0001fffc0001fffc0001fffc0001fffc0000fffc0001fff40000fffc0000fffc0000fffc00007ffc0";
 when "01100001110" => data <= 768x"0007fffe0007fffc0007fffe00077ffc0007fffe0007fffc0007fffc0007f7fc0007fffc0007fffc0007fffc00077f7c0007fff80007fffc0007fffc0007fffc0007fff80007fffc0007fff800077f7c0003fffc0007fffc0003fffc0007fffc";
 when "01100001111" => data <= 768x"0001ffff0001ffff0001ffff00017f7f0003ffff0001ffff0003ffff0001f7f70003ffff0001ffff0003fffe00017f7f0003fffe0001ffff0001fffe0001ffff0001fffe0001ffff0001fffe0001ff7f0001fffe0001ffff0001fffe0001fff7";
 when "01100010000" => data <= 768x"0000ffff0001ffff0000ffff0001ff7f0000ffff0001ffff0000ffff0001f7ff0000ffff0001ffff0000ffff00017f7f0000ffff0001ffff0000ffff0001ffff0000ffff0001ffff0000ffff00017f7f0000ffff0001ffff0000ffff0001ffff";
 when "01100010001" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff";
 when "01100010010" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff";
 when "01100010011" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0001ffff00033fff001717ff";
 when "01100010100" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f00033fff00171fff000f07ff001717ff";
 when "01100010101" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00071f7f000f0fff001717ff000f0fff001f17ff";
 when "01100010110" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff00055fff000f0fff0017177f000f0fff000f0fff000f0fff000717ff";
 when "01100010111" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00071fff00071fff001f07ff000f0fff00071f7f000f0fff00071fff00070fff00071fff";
 when "01100011000" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0000ffff00017f7f00033fff00071fff000f0fff001717ff000f0fff00071fff000f0fff00071f7f00071fff00071fff00070fff00071fff";
 when "01100011001" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff0000ffff0000ffff0003ffff00071f7f000f0fff001717ff000f0fff00071fff00070fff00071fff000f0fff00071f7f00071fff00071fff00071fff00071fff";
 when "01100011010" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff0000ffff0000ffff00055fff000f1fff0017177f000f0fff00071fff00071fff00071fff000f0fff00071fff00070fff00071f7f00071fff00071fff000f0fff00071fff";
 when "01100011011" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000177ff00033fff00171fff000f0fff0017177f00071fff00071fff00071fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff000f0fff00071fff";
 when "01100011100" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00017fff00070fff001717ff000f0fff00071f7f00033fff00071fff000f0fff00071fff00070fff00071fff00071fff00071f7f00071fff00071fff000f0fff001717ff";
 when "01100011101" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0002bfff00071fff000f0fff001717ff000f0fff00071f7f00033fff00071fff000f0fff00071fff00070fff00071fff00071fff00071f7f00071fff00071fff000f0fff001717ff";
 when "01100011110" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff00007fff00033fff00071fff00071fff000717ff00070fff00051f7f00033fff00071fff000f0fff00071fff00070fff00071fff00071fff00071f7f00071fff00071fff000f0fff001717ff";
 when "01100011111" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff00007fff00033fff00071fff00071fff00071fff00070fff00071f7f00033fff00071fff000f0fff00071fff00070fff00071fff00071fff00071f7f00071fff00071fff000f0fff001717ff";
 when "01100100000" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff00007fff00013fff00071fff00071fff00071fff00071fff00071f7f00033fff00071fff00070fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff000f0fff001717ff";
 when "01100100001" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00071fff00071fff00071fff00071fff00071f7f00033fff00071fff00071fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff000f0fff000717ff";
 when "01100100010" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00071fff00071fff00071fff00071fff00071f7f00033fff00071fff00071fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff000f0fff000717ff";
 when "01100100011" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00071fff00071fff00071fff00071fff00071f7f00033fff00071fff00071fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff000f0fff000717ff";
 when "01100100100" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00071fff00071fff00071fff00070fff00071f7f00033fff00071fff00071fff00071fff000f0fff00071fff00071fff00071f7f00071fff00071fff00070fff000717ff";
 when "01100100101" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00051fff00071fff00071fff00070fff00071f7f00033fff00071fff00071fff00071fff000f0fff00071fff00070fff00071f7f00071fff00071fff00070fff00071fff";
 when "01100100110" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00051fff00031fff00071fff00070fff00071f7f00033fff00071fff00031fff00071fff000f0fff00071fff00070fff00071f7f00071fff00071fff00070fff00071fff";
 when "01100100111" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00051fff00031fff00071fff00070fff0007177f00033fff00051fff00031fff00071fff000f0fff00071fff000f0fff00071f7f00071fff00071fff00070fff00071fff";
 when "01100101000" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff00051fff00030fff00071fff00070fff0007177f00033fff00011fff00031fff000713ff000f03ff000707ff000f0fff00071f7f000f1fff00071fff00070fff000717ff";
 when "01100101001" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000117ff00030fff000707ff00030fff0007177f00030fff00011fff00030fff000717ff000f0fff000711ff000f03ff0007077f00070fff00071fff000f0fff00071fff";
 when "01100101010" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000117ff00030fff000507ff00030fff0005177f00030fff00011fff00070fff000717ff00030fff00070dff000309ff0007077f000307ff000707ff00070fff000717ff";
 when "01100101011" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000117ff00030fff000507ff00030fff0005177f00032fff00071fff00030fff000117ff000301ff000115ff00031eff00071f7f00030fff000707ff000707ff000717ff";
 when "01100101100" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000077ff00003fff00050fff00030fff000707ff00030fff000505ff000300ff0001117700030e7f00010f7f00030fbf00031fff00031fff00071fff00070fff000707ff";
 when "01100101101" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000ffff000177ff0000ffff0000ffff0000bfff00011d7f000309ff000701ff000300ff000115ff00033cff00011dff00030cff0001177f000307ff000107ff00030fff000117ff";
 when "01100101110" => data <= 768x"0000ffff0000ffff0000ffff00017f7f0000ffff0000ffff0000efff000177ff0000efff0000dfff00008fff00011f7f00031fff00071fff000f1fff000717ff00030fff00071fff00031fff00071f7f00031fff000707ff00030fff000117ff";
 when "01100101111" => data <= 768x"0000ffff0000ffff0002ffff00037f7f0003ffff0001ffff0003ffff00017fff0001ffff0001ffff0003ffff00037f7f0003ffff00077fff00073fff00071fff000f3fff00071fff000f3fff00071f7f00073fff00071fff00030fff000717ff";
 when "01100110000" => data <= 768x"0000ffff0000ffff0004ffff00057f7f0006ffff0004ffff0006ffff0005ffff0002ffff0001ffff0003ffff00077f7f0003ffff0007ffff0007ffff00073fff000f3fff00071fff000f3fff00071f7f000f3fff00071fff000f1fff000717ff";
 when "01100110001" => data <= 768x"0000ffff0001ffff0000ffff00057f7f0006ffff0005ffff0006ffff0005ffff0002ffff0005ffff0002ffff00077f7f0003ffff0007ffff0006ffff00077fff000f3fff000f1fff000f3fff00073f7f000f3fff00175fff000f3fff001717ff";
 when "01100110010" => data <= 768x"0000ffff0001ffff0000ffff0005ff7f0006ffff0005ffff0006ffff0005ffff0002ffff0005ffff0002ffff00077f7f0003ffff0007ffff0006ffff00077fff000f3fff001f1fff000e3fff00173f7f000f3fff00177fff000e3fff001717ff";
 when "01100110011" => data <= 768x"0000ffff0001ffff0000ffff0005ff7f0006ffff0005ffff0006ffff0005ffff0002ffff0005ffff0003ffff00077f7f0003ffff0007ffff0007ffff00077fff000e3fff001f1fff000e3fff001f3f7f000e3fff001f7fff000e3fff001737ff";
 when "01100110100" => data <= 768x"0001ffff0001ffff0001ffff0005ff7f0007ffff0005ffff0007ffff0005ffff0003ffff0005ffff0003ffff00077f7f0007ffff0007ffff0007ffff000577ff000e3fff001f7fff000e3fff001f7f7f000e3fff001f7fff000e3fff001777ff";
 when "01100110101" => data <= 768x"0001ffff0001ffff0001ffff0005ff7f0007ffff0005ffff0007ffff0005ffff0003ffff0005ffff0003ffff00077f7f0007ffff0007ffff000fffff00057fff000e3fff001c7fff001e3fff001f7f7f001e3fff001c7fff000e3fff001777ff";
 when "01100110110" => data <= 768x"0003ffff0001ffff0001ffff00057f7f0007ffff0005ffff0007ffff0007ffff0003ffff0005ffff0003ffff00077f7f0007ffff0005ffff000fffff00157fff001e7fff001c7fff001e3fff001c7f7f001e7fff001c7fff000e7fff001477ff";
 when "01100110111" => data <= 768x"0003ffff0001ffff0003ffff00057f7f0007ffff0007ffff0007ffff0007ffff0003ffff0007ffff0007ffff00077f7f000fffff000fffff000fffff001d7fff001c7fff001c7fff001c7fff001c7f7f001cffff001c7fff001c7fff001c77ff";
 when "01100111000" => data <= 768x"0003ffff0003ffff0003ffff00077f7f0003ffff0005ffff0007ffff0007ffff0003ffff0005ffff0007ffff00077f7f000fffff001dffff000cffff001c7fff003c7fff001c7fff003cffff001d7f7f001cffff001c7fff001c7fff001c77ff";
 when "01100111001" => data <= 768x"0003ffff0007ffff000fffff00077f7f000fffff000fffff000fffff0007ffff000fffff001fffff001fffff001f7f7f001bffff001dffff0018ffff001c7fff00387fff001c7fff0038ffff001d7f7f0038ffff001c7fff00183fff001877ff";
 when "01100111010" => data <= 768x"0007ffff0007ffff002fffff00177f7f001fffff001fffff000fffff0017ffff0003ffff0001ffff0003ffff00117f7f00187fff00107fff00187fff00107fff0030ffff00107fff0038ffff00107f7f00003fff00507fff0008ffff00507fff";
 when "01100111011" => data <= 768x"000fffff001fffff000fffff00177f7f0009ffff001dffff000cffff001477ff000e7fff001d5fff00083fff01101f7f00001fff00107fff00007fff00107fff00007fff00107fff00003fff00501f7f00007fff00505fff00101fff00105fff";
 when "01100111100" => data <= 768x"001fffff001fffff001fffff001f7f7f001fffff001fffff001fffff001fffff0018ffff00107fff00007fff0010777f001023ff001047ff00183fff001077ff00203fff00545fff00083fff00141f7f00201fff001047ff000033ff001077ff";
 when "01100111101" => data <= 768x"003fffff001fffff001fffff001f7f7f003fffff001fffff003dffff00117ff70000ffff00005fff00007fff0010777f003867ff001047ff00380fff00101ff700203fff00501fff00001fff0010477f002073ff00107fff00003fff00001fff";
 when "01100111110" => data <= 768x"003fffff001fffff003fffff001fff7f003fffff0017ffff0003ffff00417fff0041bfff00417fff0020efff0031077f00207fff00107fff00307fff00307fff00203fff00015fff0000efff0000777f00007fff00407fff00003fff00407fff";
 when "01100111111" => data <= 768x"003fffff001fffff003fffff001fff7f003fffff0045ffff0043ffff004177ff0061ffff0041ffff0002ffff0040177f0000bfff00017fff0000ffff00007fff00023fff00417fff0040ffff00417f7f0040ffff00407fff00c0ffff0041ffff";
 when "01101000000" => data <= 768x"001fffff001fffff001fffff001f7f7f0023ffff0041ffff02e3ffff0561ffff0263ffff5745ffffffe0ffff01e07f7f00e0ffff01d5ffff00f8ffff01f17fff01ebbfff01c77fff01e3ffff0161ff7f01e3ffff01c7ffff01c3ffff01d7ffff";
 when "01101000001" => data <= 768x"0007ffff0007ffff000fffff0007ff7f0009ffff0011ffff0038ffff017077ff01b87fff75d17ffffaf83fff51703f7f00783fff007d5fff007e3fff00771fff00fbbfff00f1dfff00fbffff01f1ff7f03f9ffff01f1ffff00e1ffff0071ffff";
 when "01101000010" => data <= 768x"0000ffff0001ffff0000ffff00017f7f00023fff00071fff000e1fff001717ff00372fff55df77fffffe23ff1517177f000f03ff000fc7ff000fc7ff001757ff001f63ff001f77ff001e3fff001f3f7f007f3fff005f1fff000e3fff00151fff";
 when "01101000011" => data <= 768x"00000fff00001fff00000fff000017ff000003ff000051ff0000e0ff000171770001e27f5455f77f7fefe23f1141711f0000e03f0015717f0000e8ff000175770000e0ff0001f57f0001e3ff0001f17f0001e1ff0001f1ff0000e3ff000051ff";
 when "01101000100" => data <= 768x"0000007f0000007f0000007f0000007f00000007000001470000018300000505000007880041579c01ffff8e01551701000003800000159c000003bf0000031500000383000007c50000078b0000070500000783000007870000038f000001c7";
 when "01101000101" => data <= 768x"00000001000000010000000100000001000000000000000100000002000000170000000a0001455f0003fffe00015517000000020000001700000006000000170000000e000000070000000e0000001f0000001e0000001f0000000e00000007";
 when "01101000110" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000040500000fff00000554000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000";
 when "01101000111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000007f00000055000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01101001000" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000380000001f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01101001001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000750000003f0000000500000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "01101001010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000f80000007d0000003f000000050000000000000000000000000000000000000000000000000000000000000000";
 when "01101001011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000003e0000001f0000000fc0000007f0000003f00000017000000030000000100000000000000000000000000000000";
 when "01101001100" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000701000007c0000007c0000007f0000003f0000003fc000001fc0000007f0000001f0000000f000000070000000300000011";
 when "01101001101" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000000140000001e0000001f0000001f8000001fc000000fe0000017f0000007f0000007f0000003f8000001fc000000fe0000007f0000003f0000001f";
 when "01101001110" => data <= 768x"00000000000000000000000000000000000000000000000000000000000000000000300000007c0000007e0000007f0000003f0000005f0000003f80000017c000001fc000000fc000000fe000000770000003f0000005f0000001f8000001f0";
 when "01101001111" => data <= 768x"0000000000000000000000000000000000000000000000000000c000000170000000f8000001fc000000fc000000750000007e0000007f0000007e000000770000003f0000001f0000001f0000001f0000001f8000001fc000000f80000017c0";
 when "01101010000" => data <= 768x"00000000000000000000000000010000000180000001c0000003e000000170000001f0000001f0000000f80000017c000001f8000001fc000000f800000070000000f80000007c000000f80000007c0000007c0000007c0000007c0000007c00";
 when "01101010001" => data <= 768x"00000000000000000002000000070000000380000007c0000003c0000001d0000003e0000001f0000003f0000003f0000003f0000001d0000003e0000001c0000003e0000001c0000003e000000170000003e0000001f0000003e0000001f000";
 when "01101010010" => data <= 768x"00000000000400000002000000070000000780000007c0000003c0000001c0000003e0000007f0000003e000000370000003e0000001c0000003c0000003c0000003c0000007c0000003c0000007c0000003e0000007c0000003c0000007c000";
 when "01101010011" => data <= 768x"00000000000400000002000000070000000780000007c0000003c0000001c0000003e0000007f0000003f0000003f0000003f0000001d0000003c000000340000003c0000007c0000003c0000007c0000003e0000007c0000003e0000007c000";
 when "01101010100" => data <= 768x"00000000000000000002000000070000000780000007c0000003c0000001c0000003e0000007f0000003f0000007f0000003f0000001d0000003c0000003c0000003c0000007c0000003c000000740000003e0000007c0000003e0000007c000";
 when "01101010101" => data <= 768x"00000000000000000002000000070000000780000007c0000007c0000001c0000003e0000007f0000003e000000770000003f0000001f0000003e0000003d0000003e0000007c0000003c000000740000003e0000007c0000007e0000007c000";
 when "01101010110" => data <= 768x"00000000000000000006000000070000000f80000007c000000fc0000007c0000003e0000007e0000003e000000770000003e0000007f0000003e0000003c0000003e0000007c0000003e000000740000003e0000007c0000007e0000007c000";
 when "01101010111" => data <= 768x"00000000000000000006000000070000000f8000000fc000000fc0000007c0000003e0000005c0000003e0000007f0000007f0000007f0000003e0000003f0000003e0000007c0000003e000000740000003e0000007c0000007e0000007c000";
 when "01101011000" => data <= 768x"00000000000000000006000000070000000f8000000fc000000fc0000007c0000003e0000001c0000003e000000770000007f0000007f0000003e0000003f0000003e0000007f000000fe000001f4000000fe0000007c0000007e0000007e000";
 when "01101011001" => data <= 768x"00000000000000000006000000070000000f8000001fc000000fc0000017c0000003e0000001c0000003e000000770000007f0000007f0000007f0000007f0000007f000001ff000001be000001760000033e0000017c0000007e0000007e000";
 when "01101011010" => data <= 768x"00000000000000000002000000070000000f8000001fc000000fc0000017c0000003e0000001c0000003e0000007f0000007f0000007f0000007f8000007f000000ff000001ff000003be000007770000063e0000047c0000007e0000007e000";
 when "01101011011" => data <= 768x"00000000000000000002000000070000000f8000000fc000000fc0000007c0000003e0000001c0000003e0000007f0000007f0000007f0000007f8000007f000003ff0000077f0000063f0000047f0000083e0000007c0000007e0000007e000";
 when "01101011100" => data <= 768x"00000000000000000003000000070000000f8000000fc000000fc0000007c0000003e0000001c0000003e000000770000007f0000007f0000007f8000017f000003ff0000077f00000c3e000014770000003e0000007c0000007e0000007e000";
 when "01101011101" => data <= 768x"0000000000010000000300000007000000078000000fc000000fc0000007c0000003e0000001c0000003e000000770000007f0000007f0000007f0000017f00000fff00001d7f0000183e000010770000003e0000007c0000007e0000007c000";
 when "01101011110" => data <= 768x"0000000000010000000300000007000000078000000fc000000fc0000007c0000003e0000001c0000003e000000770000007f0000007f0000007f0000177f00001fbf00001c7f0000003e000000770000003e0000007c0000007e0000007c000";
 when "01101011111" => data <= 768x"0000000000010000000380000007000000078000000fc000000fc0000007c0000003e0000001c0000003e000000770000007f0000007f000000ff000017ff00003a3f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100000" => data <= 768x"0000000000010000000380000007000000078000000fc000000fe0000007c0000003e0000001c0000003e000000770000007f0000007f00000eff00001fff0000203f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100001" => data <= 768x"0000000000010000000380000007800000078000000fc000000fe0000007c0000003e0000001c0000003e000010770000007f0000007f00003eff0000577f0000003f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100010" => data <= 768x"0000000000010000000380000007800000078000000fc000000fe0000007c0000003e0000001c0000003e000000770000007f0000147f00003eff0000177f0000003f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100011" => data <= 768x"00000000000100000003800000070000000780000007c000000fe0000007c0000003e0000001c0000003e000000770000007f0000547f00007fff0000077f0000003f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100100" => data <= 768x"00000000000100000003800000070000000780000007c000000fe0000007c0000003e0000001c0000003e000000770000007f000054ff00003fff0000057f0000003f0000007f0000003e000000770000003e0000007c0000003e0000007c000";
 when "01101100101" => data <= 768x"0000000000010000000380000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000000ff000054ff00003fff8000057f0000003f0000007f0000003e0000007f0000003e0000007c0000003e0000007c000";
 when "01101100110" => data <= 768x"0000000000010000000380000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000000ff000054ff00000fff8000057f0000003f0000007f0000003e0000007f0000003e0000007c0000003e0000007c000";
 when "01101100111" => data <= 768x"0000000000010000000180000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000000ff000074ff00000fff8000057f0000003f0000007f0000003f000000771000003e0000007c0000003e0000007f000";
 when "01101101000" => data <= 768x"0000000000010000000180000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000020ff000055ff00000fff8000057f0000003f0000007f0000003f000000771000003e0000007c0000003e0000007f000";
 when "01101101001" => data <= 768x"0000000000010000000180000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000020ff000055ff00000fff8000057f0000003f0000007f0000003f000000771000003e0000007c0000003e0000007f000";
 when "01101101010" => data <= 768x"0000000000010000000180000007c000000780000007c000000fe0000007c0000003e0000001e0000003e00000077000020ff000055ff00000fff8000057f0000003f0000007f0000003f000000771000003e0000007c0000003e0000007f000";
 when "01101101011" => data <= 768x"0000000000010000000180000007c00000078000000fc000000fe0000007c0000003e0000001e0000003e00000077000020ff000074ff00000fff8000057f0000003f0000007f0000003f000000771000003e0000007e0000003e0000007f000";
 when "01101101100" => data <= 768x"0000000000010000000380000007c0000007c000000fc000000fe0000007c0000003e0000001e0000003e00000077000000ff000075ff00002fff8000057f0000003f0000007f0000003f000000770000003e0000007f0000007e0000007f000";
 when "01101101101" => data <= 768x"0000000000010000000380000007c000000fc000000fc000000fe0000007c0000003e0000005e0000007e00001077000030ff000055ff00002fff8000057f0000003f8000007f0000007f000000770000007e0000007f0000007e00000077000";
 when "01101101110" => data <= 768x"000000000001c0000003c00000074000000fc0000007c000000fe0000007e0000003e0000005f0000007e00001077000030ff000055ff00002fff8000057f0000003f8000007f0000007f800000770000007f0000007f0000007e00000077000";
 when "01101101111" => data <= 768x"000000000001c0000007c000000740000007e0000007c0000007e0000007f0000003e0000005f0000007f00003077000030ff800055ff00000fff0000057f0000003f0000007f0000007f800000770000007f0000007f000000fe0000007f000";
 when "01101110000" => data <= 768x"0000000000004000000fe0000007d0000007e0000007c0000007e0000007f0000003e0000007f0000307f00007077000030ff800055ff40002fff8000057f0000003f8000007dc000007e800000771000007f8000007f000000fe0000007f000";
 when "01101110001" => data <= 768x"0000000000045000000ef0000007f0000003e0000007c0000007e000000770000003e0000107f000038ff00007077000030ff800055ff40002fff8000077f0000003f8000007dc000007ec00000775000007e8000007f000000ff0000017f000";
 when "01101110010" => data <= 768x"0000000000041000000e30000007f0000003e0000007e0000007e0000107f0000207e0000507f000038ff80007077000030ff000075ff00000fff0000077f0000003f8000007f4000003e600000777000007f2000007f000000ff8000007f000";
 when "01101110011" => data <= 768x"0000000000040000000730000007f0000003f0000007f0000007e0000107f0000307e0000507d000038ff00007077000030ff000075ff00000fff0000077f0000003fc000007c5000003e380000771000007f0000007f000000ff8000007f000";
 when "01101110100" => data <= 768x"0000000000040000000780000007f0000003f0000007f0000007e0000107f0000307e0000747c000038fe000071ff000031ff000055ff00000fff000007f70000027fe000007c7000003e380000771000007f0000007f000000ff8000007f000";
 when "01101110101" => data <= 768x"0000000000050000000780000007f0000003f0000007f0000007e0000107f0000387c0000547c000038fe000071ff000033ff000055ff00000fff000007f7000003ffe000017c7c00003e1c0000771000007f0000007f000000ff8000007f000";
 when "01101110110" => data <= 768x"0000000000050000000380000007f0000003f0000007f0000007e0000107f0000387c0000547c000038fe000031f7000031ff000055ff00000fff000007ff500003fff800017c5c00003e080000770000007f0000007f000000ff8000007f000";
 when "01101110111" => data <= 768x"0000000000050000000380000007f0000003f0000107f0000007e0000107f0000287c0000547c0000387e0000307f000038ff000055ff00000fff000007ff500001fff80000fc5c0000fe000000770000007f0000007f000000ff8000017f000";
 when "01101111000" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000287c00001c7c000038fe0000307f000038ff000055ff00000fff800007ff5400007efe00007c5400003e000000770000007f0000007f000000ff8000017f000";
 when "01101111001" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000187c00001c7c000038fe00003077000038ff000054ff00000fff800007ff540000fffc00007c0000003e000000771000007e0000007f000000ff0000017f000";
 when "01101111010" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000287c0000107c000038fe0000307f000038ff000055ff00000fff800007ff540000fef800007c0000003e000000771000007e0000007f000000ff0000017f000";
 when "01101111011" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000007c0000147c000038fe00003c7f000038ff000055ff00000fff800007fd540000fef800017c0000007e000001771000007e0000007f000000ff0000017f000";
 when "01101111100" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000307c0000547c000038fe0000347f000030ff000055ff00000fff800007fd540000fefa0001fc1000007e00000077000000fe0000007f000000ff000001ff000";
 when "01101111101" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000387c00005c7c000038fe0000307f000030ff000055ff00000fff800007fd550000fefe0001fc1000007e0000007e000000fe0000007f000000ff000001ff000";
 when "01101111110" => data <= 768x"0000000000010000000380000007f0000003f0000007f0000007f0000107f0000387c0000547c000038fe0000707f000030ff000075ff04000fff800005fd500000fefe00007c1000007e0000007e000000fe0000007f000000ff000001ff000";
 when "01101111111" => data <= 768x"0000000000050000000380000007f0000003f0000107f0000007f0000107f0000307c0000507c000038fe0000707f000030ff000075ff04000fff8c0005fd540000fefe00007c1400007e0000007e100000fe0000007f000000ff0000017f000";
 when "01110000000" => data <= 768x"00000000000500000007a0000107f0000003f0000007f0000007e0000107f0000307c0000507c000038fe00007077000030ff000075ff04000fff8c0007fd540000fefe00007c1400007e0000007e100000fe0000007f000000ff0000017f000";
 when "01110000001" => data <= 768x"00000000000400000007a0000107f0000003f0000007f0000007e0000107f0000307c0000707c000038fe000031ff000030ff000055ff04000fff8e00077d540000fefe00007c1400007e0000007e100000fe0000007f000000ff000001ff000";
 when "01110000010" => data <= 768x"00000000000400000007b000000770000003f0000007f0000007e0000107f0000387e0000507c000038fe000011f7040031ff0e005dff04000fff0400077d740000fefa00007c0000007e00000077000000fe0000007f000000ff000001ff000";
 when "01110000011" => data <= 768x"0000000000040000000630000007f0000003e0000107f0000087e0000147e0000387e00001c7c14001cfe0c0011f71c0038ff1c001dff04000fffa800077df40000fea000007c0000007e00000077000000fe0000007f000000ff000001ff000";
 when "01110000100" => data <= 768x"0000000000040000000e3000000770000003e0000147c10000e7e0000157c10000e7e38000c7c5c000cff380015f710000eff300007ff740003ffe000037dc00000ff8000007c0000007e00000077000000fe0000007f000000ff000001ff000";
 when "01110000101" => data <= 768x"0000000000040000000e20000017f1000027e0000057c4000077e6000177d7000077e7000077c700008ff600015f7700003ffe00007ffc00003ffc000017f400000ff0000007c0000007e000000770000007e0000007f000000ff000001ff000";
 when "01110000110" => data <= 768x"0000000000000000000e70000017f000003fea000057cc00003fee000077df000037ee000057c400006ffe00017ff400003ffc00001ffc00001ff8000007f000000ff0000007c0000007e000000770000007e0000007f000000ff000001ff000";
 when "01110000111" => data <= 768x"0000000000000000000c30000017f400003ffa000057dc00003fee000077d4000037ec000057c400003fec00013f7c00003ff800001ffc00000ff8000007f000000ff0000007d0000007e000000770000007e0000007f000000ff000001ff000";
 when "01110001000" => data <= 768x"000000000050040000083200005f7500003ffe00007fdf00007ffe000077fc00003fee000057e400003fec0001377c00003ffc00001ffc00001ff8000017f000000fe0000007f0000007e000000740000007e0000007f000000ff0000017f000";
 when "01110001001" => data <= 768x"002002000054550000783e00017d7f0000ffff00017fff0000fffe000077f700007ffe000057f5000067ee0000777c00003ffc00001ffc00003ff8000017fc00000ff0000017f000000ff000000770000007e0000007c000000fe0000017f000";
 when "01110001010" => data <= 768x"00f82f8001f5554001f83f8001fd770003ffff0001ffff0000ffff8001f7f70001ffff8001fff70000ffee000077f500003ffe00007ffc00003ffc000037fc00003ff8000017f000000ff00000177000000ff0000007f000000fe0000007f000";
 when "01110001011" => data <= 768x"03fa238005d5554006fe7f80057f775003fe3f8005fd7f4003ffffc007f77fd003ffffc005ffff4003ffff8001f7f70000efee000077ff0000fffe00007ffc00003ffe00007ffc00003ffc00001ff000000ff000001ff000000ff8000017f000";
 when "01110001100" => data <= 768x"03fe2ec005fd55c003fe0fc01755574007fe3f8007fc5fd00ffeffe017fffff007ffffe017ffffc00fffff80077f774003ffff8001dff70000efff0001f7f70000fffe00007ffc00007ffe00007f7400003ffc00001ff000000ff800001ff000";
 when "01110001101" => data <= 768x"1fba0fe01dd557500ffe2fe0177d57741bfe2ff817fd5ff50ffe3ffa57fd7ff43ffffff857ffffd00fffffe0177f7fd00fffffe007dff7c003efffc001d7f74001efff0001dff70000ffff00017f7f0000fffe00007ffc00003ffe00001ff400";
 when "01110001110" => data <= 768x"23bbaff257d557f42ffbaffc577757753ffa3ffe5ffd5ffc7ffe3ffc7fff77f43ffe3fe85ffd5ff41ffffff85f7ffff03ffffff05fffffd00fffffe007d7f77003efffc001dff74003efff80015f770001ffff0001ffff0000fffe00007ff700";
 when "01110001111" => data <= 768x"1ffbbfa35ff55f57bff8bfee57757f55fffa3ffa7ff55fd5fffefffa77f557f53ffebffa7ffd5ffc3ff83ffc7f7d7f743ffffff85ffffff43ffffff817fffff01ffffff01ffffff00fffffe007df77c103dfff8007dff78003ffff80017ff700";
 when "01110010000" => data <= 768x"a3fbfff857fdfff53ffefff857fd7f753ffe3ffa7ffd5ffdfffebffe7fff57f5fffebffe7ffd5ffcffff9ffc7f7d5f7d3fffbffe5ffffffd3ffffffc5fff77f43ffffff81ffffff40fffffe0155f77503e1ff2381f1ff1f00f9ffbf817dff7f0";
 when "01110010001" => data <= 768x"ffff3ffa7fff5ffdffff3ffe7f7f1f7dffff3fff7fff5ffdffffbffe77ff7ff77fffffff7ffd7fffffffffff7f7f7f7f7ffffffe7fffffff7fffbffe77f77ff73ffffffe5ffffffc0ffffffc577f777403fffff0055ff550000ff0001017f110";
 when "01110010010" => data <= 768x"afbfbfff577f5ffdafffbfff57ff5f7f3fffbfff7fff7fffffffffff77f7f7ffffffffff7fffffffffffffff7f7f7f7fffffffff7fff7fffffffffff7ff77fff3ffe3fff5ffd5fff3ffebfff5f7f7fff1ffffffe17fffffc03fffff8011ff550";
 when "01110010011" => data <= 768x"ffffffff7fffffffffffffff7f7f7f7fffffffffffffffffffffffff77f7ffffffffffffffffffffffffffff7f777f7fffffffffffffffffffffffffffffffffffffffff7fffffff3fffffff7f7f7f7f3fff3fff5ffffffd3ffffffe577ff7f5";
 when "01110010100" => data <= 768x"fffffffbfffffff5ffffffff7f7f7f7ffffffffffffffffffffffffffffffff7ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7fffffffffffffffffffffffff5ffffff7";
 when "01110010101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffff7fffdfff";
 when "01110010110" => data <= 768x"fffffffffffdffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110010111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7dfffffffffffffffdfffffffffffffff7ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011000" => data <= 768x"ffffffffffffffdfffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011011" => data <= 768x"ffffffffffffffffffffffff7f7f7f77ffffffff7fffffffffffffff7ffffff7ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffff7fffffff";
 when "01110011101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffff5fffffffffffffffdffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011110" => data <= 768x"fffffffbfffffff5fffffffe7f7f7f7dffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffff7ffff7ffffffffffffffffffffffffffff7f7f7fffffffffffffffffffffffffffffffff";
 when "01110011111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f777f7ffffffffffffffffffffffffff7ffffff";
 when "01110100000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffff77ffffffffffffffffffffffffffffff7f5f7f7fffbfffffff5fffffffafffff77d7ffffffffffff7fdfffffffffffff7f777f7fffffffff5ff7ffffbfffffff57f5ffff";
 when "01110100001" => data <= 768x"fbffffff55d7ffffffffffff5f777f7fbfffffff5fd7ffffafefffff57d7ffff2fffffff57d7ffff0fffffff17d77f7f0fffffff5fffffff3fffffff5fffffff3fffffff5ff7ffff3fffffff7ff77f7f3fe3ffff1fd5ffff0703ffff0511ffff";
 when "01110100010" => data <= 768x"022fffff1557ffff38afffff1d577f7f1e3fffff1d5fffff1eafffff1f57ffff0fafffff1fd7ffff0f8bffff1f557f7f0f83ffff17d5ffff1fc3ffff17d5ffff1fe3ffff1fc5ffff3fe3ffff7f577f7f3fe3ffff1fc5ffff0703ffff1505ffff";
 when "01110100011" => data <= 768x"000bbfff40555fff300bffff7d177f7f3e07ffff1c17ffff1e0fffff1f17ffff1f83ffff1f15ffff3f83ffff3f157f7f3f8bffff17d7ffff2fcfffff17d7ffff1fefffff1fd7ffff3fefffff7ff77f7f3fe3ffff1fc5ffff0703ffff05157fff";
 when "01110100100" => data <= 768x"0003ffff0005ffff2003ffff7c157f7f3c0bffff1c15ffff3e0fffff1717ffff3f8fffff7f57ffff7f8fffff77577f7fffbfffff17d7ffff2fefffff17d7ffff1fefffff1fd7ffff3fe7ffff7ff77f7f3fe3ffff1fd5ffff0700ffff05117fff";
 when "01110100101" => data <= 768x"0023fffb0055fff520afffff75577f773c3fffff1d57ffff3ebfffff1757ffff3fbfffff7f57ffffff8ffffff7577f7fd78fffff57d7ffff2fcfffff07d7ffff0fffffff1fd7ffff3fefffff3ff77f7f3fe3ffff1fc57fff0700ffff05117fff";
 when "01110100110" => data <= 768x"000fffff0157ffff000fffff75177f7f380fffff1c1fffff3c0fffff1f17fff73f8fffff7f17ffffff8ffffff7177f7ff78fffff57d7ffff2fcfffff07d7ffff0febffff1fd5ffff1febffff3f557f7f3fe3ffff1fc5ffff0703ffff0515ffff";
 when "01110100111" => data <= 768x"003fffff005ffdfd003fffff751f7f7f782fffff5d57ffff3e0fffff1f57fff73f8fffff7f57ffffff8fffff77577f7fffafffff57d7ffff278fffff07d7ffff0fefffff1fd7ffff1fefffff3f77ff7f3fefffff1fd5ffff070fffff0515ffff";
 when "01110101000" => data <= 768x"002bffff1555ffff000fffff75177f7f780fffff5c57ffff3c0fffff1f17ffff3f0fffff7f57ffff7fbfffff775f7f7f7fbfffff57dfffffa7ffffff07dfffff0fffffff1fdfffff1fefffff3f777f7f3febffff1fd5ffff0703ffff0517ffff";
 when "01110101001" => data <= 768x"003fffff0057ffff003fffff71577f7f783fffff5d5fffff3cffffff1f77ffff3fbfffff7f5fffff7fbfffff77577f7f7fbfffff77d7ffff678fffff07d7ffff0fe3ffff1fd5ffff3febffff3f577f7f3fefffff5fd7ffff0f8fffff0557ffff";
 when "01110101010" => data <= 768x"00ffffff015fffff00ffffff71577f7f783fffff5c57ffff3c2fffff1f57ffff3fabffff7f57ffff7f8fffff77177f7f7f8fffff7757ffff6f8fffff17d7ffff0fffffff1fd7ffff3fffffff3f777f7f3fffffff5fd7ffff0fcfffff0557ffff";
 when "01110101011" => data <= 768x"0003ffff0055ffff000fffff71177f7f780fffff5d57ffff3c0fffff1f57ffff3fafffff7f57ffff7f8fffff77177f7f77afffff77d7ffff77bfffff17dfffff0fffffff1fdfffff1fefffff1f577f7f3fefffff5fd7ffff0fcbffff0515ffff";
 when "01110101100" => data <= 768x"003fffff045fffff000fffff71577f7f383fffff5d5fffff3c3fffff1f57ffff3fbfffff7f5fffff7fffffff7f7f7f7f7fbfffff77dfffff7fffffff17dfffff0fffffff1fdfffff1fffffff1f777f7f3fffffff5fd7ffff0fcfffff0515fff7";
 when "01110101101" => data <= 768x"00bbffff05557fff00feffff75557f7f3bfbffff5d557fff3efeffff1f557fff3ffbffff7fd5ffff7faaffff77557f7f7fbbffff77d5ffff7f8fffff17d7ffff0fffffff1fd5ffff1fe3ffff1fd57f7f3fe3ffff5fc5ffff0fc2ffff05157fff";
 when "01110101110" => data <= 768x"0203ffff5555ffff0a8bffff75577f7f3f0fffff5d57ffff3e8fffff1f57ffff3f0fffff5f57ffff3f8fffff7717ff7f7f8fffff7757ffff778fffff17d7ffff0fc3ffff1fd5ffff1fe0ffff1f557f7f3fe03fff5fd55fff0fe80fff055517f7";
 when "01110101111" => data <= 768x"000fffff1557ffff000fffff55177f7f3e0fffff1c17ffff3e0fffff1517ffff3f0fffff5f17ffff3f8fffff7f177f7f7f83ffff77557fff7f80fffe17d57fff0fc03fff1fc55fff1fe03fff1f6117ff3fe03fff5fe157ff0fc00fff051157f5";
 when "01110110000" => data <= 768x"000fffff0017ffff000fffff55177f7f3c0bffff1c15fffd3c0affff15157ff53f00fffb5f155ff53f803ffa7f0117757f802ffb770055f57f800ffe17c117ff0fc02bff1fc055ff1fe00fff1f61577f3fe02bff7fe155fd0fc02fe805115571";
 when "01110110001" => data <= 768x"00003efa00005d5d00003efa140015753c000bfa1c0015751e000bf8150015f53f0003f25f0005f53f8003f07f1117717f8003f0778505f17f8003f817d515f50fc203fe1fc515fd1fe003fe1fd515ff3fe003ff7fe015fd0fc000e805001171";
 when "01110110010" => data <= 768x"000000000000054400000008100001703e0000781c0005781e0000781f0001703f0001f01f0001f03f8001f07f0101707f8001f0770005f07f8001f817c101fc0fc003fe1fc001ff1fe003fe1fc0017f3fe003fe7fc001fc0fc000e005000140";
 when "01110110011" => data <= 768x"000000000000000400000008140000713e0000781c0000701e0000781f0001703f0001f81f0001fc3f8001fc7f0001747b8001fe778001f46f8003f817c001fc0fc003fe1fc001fc1fe003fe1fc0017f3fe003fe7fc001fc0fc000e005000140";
 when "01110110100" => data <= 768x"000000000000000000000008140000703e0000701c0000701e0000781f0001741f0001fe1f0001c73f8001e7770001577b8003f2778001f44f8003f817c0017c0fc003fe1fc007fc1fe003fe1f40077f3fe003fe7fc005fc0fc001e005000140";
 when "01110110101" => data <= 768x"000000000000000000000008140000701e0000701f0000700e0000781f0001f41f8001fe1fc001ff3f8001ef7fc001517b8003f057c001d00fc003f817c001700fc003fc1fc007fc1fe003fe1fc0077f3fe003fe5fc007f40fc001e005000140";
 when "01110110110" => data <= 768x"000000000000000400000008150000700f000070070000700f0000f8170001f01f8003fc1fc001ff3fc003ff77c001557fc003f655c001f40bc003f817c003f007e003f807c007fc0fe007fc1f70077c3fe007fe1ff007f40fe000e007000140";
 when "01110110111" => data <= 768x"00000000000000100000002007000170038000f007c001f0078000f0074001f00fc003f81fc007fc3fe003fe3f4103773be003f257c007f007e003f805f007f003f003f807f007fc0ff007fc1f70077c3ff007fc17f007f407e001e001400140";
 when "01110111000" => data <= 768x"0000000004000040010000c0014001c003e003e001c001c003c001e007c003700fe003f81ff007fc1ff007f81571077d3bf007fc117007d403f007e007f007f003f007f807f007fc0ff807fc17f0077d1ff807f817fc07f003f803c001500140";
 when "01110111001" => data <= 768x"000000000040010000e001000041070000f0078001f007c003e003e0074003700fe003381f70071c3ef80f9c75f007d431f0078611f0074000f007e001f0077001f007f805f007fc07f807fe17f007ff1ff807fe1ff007fd3ff803fc17f00370";
 when "01110111010" => data <= 768x"002000000010040000300c000070050000f00f0001dc1fc003f80ff817f007ff3fe003ff7f70075ffe700f0375700701e0f80f0040f0070000f00f800070074000f007e001f007f403f007fe0770077f0ff007ff1ff007ff7ff00fff7ff007ff";
 when "01110111011" => data <= 768x"000000000004100000081000001c100000381e00007c1f0000fc3f8007fc3ff53ff83fff7ff017ffffe007ff7d710715f8f22f0050f44f0000fe3f000174770000fe3f0001fc1f0001e007e0037107f103e007fe07f007ff1fe007ff77f007ff";
 when "01110111100" => data <= 768x"00000000000100000002000000157000001c3000007c1d0000fc3f0001fc770003fe3fe017fc5ffd3ff80fff7f70077ffff18ffffff11f7ffff98ffff5f75f5181fbbf8001f75f0001fe7f80017017c003e007f007e007fc0fe007fe1ff007ff";
 when "01110111101" => data <= 768x"00000000000100000002000000154000000e2000007c1d0000fc3f0001fc770001fe7f8001fc5fc007f81ff81770177d3ff91fff7ff11ffffff99fff7f77dff5bffbbfbe75f75f15e1fe7f800170174003e007f007f007fc07e007fc17f007f4";
 when "01110111110" => data <= 768x"00000000000100000002000000154000000e2000007c1c0000fc3f0001fc770000fe3f0001fc5f0001f81f80017017c003f81fe007fd1ff00ff9bff01fff7ff01ffbbff81dff5fdc3bfe7fc007f4574003e807e007f047f407e007fc17f007fc";
 when "01110111111" => data <= 768x"00000000000000000002000000154000001e2000007c1c0000fc3f0001f4770000fe3f0001fc5f0000f80f800170070003f00f8001f11fc003fb8fc003f7ffc003ffbfc007fd7fc003fe7fc0037517c003e20ff007f107fc07e00ffc07f007fc";
 when "01111000000" => data <= 768x"00000000000000000002000000154000001e2000007c1c0000fc3f0001f4770000fe3f0001fc5f0001f80f8001f0070001f00f8001f11fc003fb8f8001f7ffc001fbbf8001f75f0001fc3f800170174003e007f007f007fc07e00ffc07f007fc";
 when "01111000001" => data <= 768x"00000000000100000002000000154000001e2000007c1c0000fc3f0001f4770000fe3f0001fc5f0001f80f8001f0070001f00f8001f11fc003fb8f8001f7ffc003fbbf8001f75fc003fc3fc0017017c003e007f007f007fc07f00ffc07f007fc";
 when "01111000010" => data <= 768x"00000000000100000002000000155000001e3000007d1c0000fc3f0001f47f0000fe3f8001fc5f0001f80f8001f0070003f00f8001f11fc003fb9fc003f7ffc003fbbfc007f75fc003fc3fe00770174003e007f007f007fc07f00ffc077007f4";
 when "01111000011" => data <= 768x"000000000004000000060000001d5100003e3800007d1d0000fc3f0001fc7f0000fe3f8001fc5f0001f81f8001f0178003f18f8001f19fc003fb9fc007ff7fc003fbbfe007ff7fc007fc3fe007f0175003f00fe007f007f003f00ff807f017fc";
 when "01111000100" => data <= 768x"00000000001440000018000000744700003e2e00007c1f0000fc3f0001fc7f0001fe3f8001fc5f0001f81f800175170003f99f8001fd9fc003fb9fc003f77fc003fbbfe007ff7fc003fc3fe007f0174003f00fe005f00ff003f00ff807f017fc";
 when "01111000101" => data <= 768x"0028000000144000003800000074410000382300007c1d0000fc3f00017c770000fe3f0001fc5f0000f83f8001f5170001f9bf8001fddfc003ffff8001f57fc003ffffc003ff7fc003fc3fc0037017c003f80fe001f01ff003f80ff8077017fc";
 when "01111000110" => data <= 768x"0010000000544000003000800074414000382100007c1d0000fc3e0000747f0000fe3f0000fc7f0000fc3f00017d3f0000ffbf0001fd5f0001ffff8001ff770001ffff8001ff7fc001fc3f8001f11f4001f80fe001f41ff003f80ff803f01ffc";
 when "01111000111" => data <= 768x"0010000000544000003000800074414000382100007c1d00007c3e0000747f0000fe3f00007c7f0000fc3f00007d7f0000ffbf0000fd5f0000ffff0001f7770001feff8001ff7f0000fc3f8001f91f0001f81fe001f01ff003f80ff803f01ff4";
 when "01111001000" => data <= 768x"0010000000544000003000800074414000382100007c1d00007e3e0000747f0000fe3e00007c7f0000fe3e00007d7f0000ffbf00007dff0000ffff00017f770000feff0001fc7f0000fc3f00017d1f0001f81fe001f01ff003f80ff801f81ff0";
 when "01111001001" => data <= 768x"0010000000544000003000800074414000382100007c5d00007e3e0000767f00007e3e00007c7f00007e7e00007d7f00007fbe00007dff0000fffe00007f770000feff00007c7f0000fe3e00007c7f0000f83fe001f01ff003f80ff801fc1ff0";
 when "01111001010" => data <= 768x"0010000000544000007000800074414000382100007c5d00007e3e0000767f00007e7e00007c7f00007e7e00007d7f00007ffe00007fff00007ffe00007f7f00007e7e00007c7f00007e3e0000747f0000f83fe001fc1ff003f81ff801fc1ff1";
 when "01111001011" => data <= 768x"0010000000544000007000800074414000382100007c5d00007e3e0000767f00007e7e00007c7f00007e7e00007d7f00007ffe00007ffc00007ffe00007f7700007efe00007c7e00007e7e0000747f0000fa3fa001fc5ff001f81ff801fc1ff0";
 when "01111001100" => data <= 768x"0010000000544000007000800174414000382000007c5d00007e3e0000767f0000fe3e00007c7f0000fe7e00007f7f00007ffe00007fff00007ffe0000777700007ffe00007f7e00007e7e00007e7f0000fe3f8001f45fd001f80ff001f01ff0";
 when "01111001101" => data <= 768x"0090000001500040007020000174014000782080007c1d00007e3f000074770000fe3f00007c7f0000fe3f00007f7f0000ffff00007fff0000fffe00007f7700007ffe00007f7f00007e7e00007c7f0000fe7e0001f45f4001f81fe001701ff0";
 when "01111001110" => data <= 768x"00f800000070100000380000017c107000382060007c154000fe3f8000773f0000fe3f8000fc7f0000fe3f80017f7f0000ff7f0001ffff0000ffff0001fff70000fffe0001fdff0000fefe00017d7f0000fcfe0001fc7d0003f8fe0001505f50";
 when "01111001111" => data <= 768x"003800000054040000fe080000741110007e0838007f041400ff0f2001ff1f5000ff1fc001ff1fc001fe3fc001ff3fc003fe3f8001ff5f0003ffff80017fff0003ffff0001ffff0003fffe0003757f0003fbfe0005f1fc0003f9fe0001517400";
 when "01111010000" => data <= 768x"003e0000005f0000003e0000017f050000ff820201ffc40500ffc20e01f7c75501ff87e801ff17d003fe1fe007fc1fc003fc3fe007fd7fc007ffffc0077fffc00fffff8007ffff000fffff0017777f000feffe0005d7fc0000e7fe0000077c00";
 when "01111010001" => data <= 768x"001fc000005fc000007f8000017fc10000ffe00001ffd10003ffe000037f710103ffe18307ffc1d50ffe03f217fc17740ffc1ff01ffd7ff01fffffe01ff777f03fffffe05fffffc03fffff80177f7f0003bffe00015ffc00001ffe000017fc00";
 when "01111010010" => data <= 768x"003ff000007fd00000ffe00001ff700003fff80007fffc4007fff80017f7fc411ffff8001ffff0403ff8a0e0777c01713ff803fb7ffd17fdfffffffc77fff7f07ffffff05ffffff00fffffe007ff7fc003ffff80017fff00007ffe00001ffc00";
 when "01111010011" => data <= 768x"007ffe0001fffc0001fff80007fffc0007fffe001ffffc001ffffe005fffff103ffffe007ffdfc10fff87e207f711410fffc00207f7c007cffff01fc5fff57fd1ffffffe07fffffd07fffff807ff7f7003ffffe001ffffc000ffff00007ffd00";
 when "01111010100" => data <= 768x"003fff0001ffff0003ffff8007ffff010fffff001fffff003fffff807ff7ff00ffbfff80ff7c7f00fffc7f887f7c3f113ffc3f005ffc1c100ffe082017f700500fff80f807ffd5fc07fffff807ff7f7503fffff201ffffc401ffff80017ffd10";
 when "01111010101" => data <= 768x"00ffff8005ffffc00fffffe01f7f7f703fffffe07fdfffd0ffffffc077f7ffc03fffffe05fff5fc01ffe3fc01f7c1fc01ff83f801ffc7f040ff87f0817f47f100ffc382007fc00400fff008007ffd75007fffff007fffff503ffffeb01fff755";
 when "01111010110" => data <= 768x"03ffffe01ffffff03fffffe0177f7f703ffffff01ffffff00ffffff81ff7f7f00ffffff81fffdff01ff81fe01f701f711ff01fe01ff05fc01fe3ffc01ff7f7c01ff3ff801ff1fd100ff8f8001f7c11400ffe020007ff55400fffff8007f77741";
 when "01111010111" => data <= 768x"0fffffb807ffffdc0ffffff8077f7f7c03fffff807fff7fc0ffffff807fffffc0ffbfff81ff07ffc1fe07ffc1f417f7d3f9c3ff81fdc1ff03f9e3fe017d77fc03f9fffc01fdfffc03fefff001f75fd003ff0b0001ffc05001fff80001577d500";
 when "01111011000" => data <= 768x"03fffe00007fff4400ffffe2017f7f7703fffffe07dfffff0ffffffe1ff07ffd1fce3ffe1fdc1ffc3fbe1efc3f7d1f7c3f783ffc7f7c7ffc3f7cfff87f777ff03f3ffff07f3fffd07f9fffc07fd77f003fe3fe0005f1540000f80000007d5400";
 when "01111011001" => data <= 768x"003ffe00007fff0000ffff80017f7fd107fffff007f57ff10fefbffb175f57fd3f3fefff1f7dd7ff3efaeffe7d75577d7efa2ffe7dfd5ffcfefffffc7577ff7cfefffff85d7ffdf02f3fffe0171f7fd1038fff8001c7fd0000e0e80000710100";
 when "01111011010" => data <= 768x"003ffe00017fff0003ffff80077f7fc10fffffe01fdfdfd01fffffe0177ff7f13ffffff87dfd77fdfdffffff7df7777ffbfffffe7dfd5ffc7dfffff85dff77f10dfffff00dfffff00effffe0077f7fc0033fff800157fd0000c2e80000510000";
 when "01111011011" => data <= 768x"01fff80005fffc000ffffe001f7f7f013fffff805fffffc07fffff8077f7ffd1ffffffe07fffdfd0ffffffe87f7fff753ffffff85ffffff03fffffe017f777d11fffff801dffff000ffffe00057ffd01033ff800055554000080000011511110";
 when "01111011100" => data <= 768x"3ffffa007ffffd40fffffe007f7f7f11ffffff00ffffff40ffffff80ffffff51ffffff80ffffff50ffffff807f7f7f51ffffff80ffffff44fffffe007ffff7513ffffe005ffffd401ffff800177f55110fffa000155554000008000011151110";
 when "01111011101" => data <= 768x"fffff800fffffd40fffffe007f7f7d11fffffe00fffffd40fffffe00ffff7d11fffffe00fffffd40fffffe007f7f7d11fffffa00fffff540fffff800fffff511ffffe0007fff54403fff80001775511102aa0000455544000000000011111110";
 when "01111011110" => data <= 768x"ffffe000ffffd400ffffe0007f7f5501ffffe000ffffd401ffffe001ffffd111ffffe000ffffd400ffffe0007f7f5101ffff8000ffff5400fffe00007ff511103fe2000055554000000000001511110000000000040400010000000111111001";
 when "01111011111" => data <= 768x"fffe0000fffd4000fffe00007f7f1101fffe0000fffd4005fffe0003f7fd1113fffa0001fff54000fff800007fd51101ffa000015554000008000000151110010000000044400001000000011111000100000003000000070000000311100007";
 when "01111100000" => data <= 768x"fff00000fff40000fff800007f710100fff00000fff40015ffe0000fffd11007ffa00003ff500005fe00000355110007000000034400000500000003111010030000000300000007000000070101000700000007000000070000000f00000017";
 when "01111100001" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40014ff80003eff51101ffe00001f554000070000000f1111001f0000000f040000070000000f111000070000000f0000001f0000000f0101001f0000001f0000001f0000001f0000001f";
 when "01111100010" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc40050ff80007cff511174fe00003e5540001f0000000f1111001f0000001f0400001d0000000f1110001d0000001f0000001f0000001f0101001f0000003f0000001f0000003f00000017";
 when "01111100011" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40050ff8000f8ff51007cfe00003e5540001c0000003f1111013f0000003f0400001d0000001c1110001d0000003e0000007c0000003e0101003f0000003f0000007f0000003f0000007f";
 when "01111100100" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc40140ff8001e0ff5111f0fe0000f85540007c0000007e1111007f000000ff0400007d000000791110007d000000f8000000fc0000007c0101007c0000007e0000007f0000007f0000007f";
 when "01111100101" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40540ff8003e0ff5111f0fe0001f055400070000000f81111017c000000fe04000057000000fb111001f1000001f8000001fc000000f80101017c000000fc000001fc000000fe000001ff";
 when "01111100110" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40540ff8003c0ff5113c0fe0003e0554001f0000000f011110170000001f8040001fc000000fe11100177000003f0000005f0000001f8010101f1000003f8000001fc000003fc000001fc";
 when "01111100111" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40500ff800780ff5107c0fe0003e0554001e0000001e011110170000003f0040001f0000001f8111001f0000003f8000005f0000001e001010170000003f0000007f0000007f8000007fc";
 when "01111101000" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40500ff800780ff5107c0fe0003e0554001c0000001e011110170000003e0040001c0000001e011101170000003e0000001d0000003e001010370000003f0000007f0000007f8000007f4";
 when "01111101001" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40500ff800780ff5107c0fe0003c0554001c0000003e011110750000003e0040001c0000003e011101140000003e0000005c0000003e001010770000003f0000007f0000007f8000007f0";
 when "01111101010" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40500ff800f80ff5107c0fe0003c0554001c0000003c011110740000003e0040001c0000003e0111013c0000003c0000007c0000003e0010107e0000007e0000007f000000ff8000007f0";
 when "01111101011" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41500ff800f80ff510700fe000380554001c0000003c011110740000003e004000740000003e011100760000003e0000007c0000007c0010107c0000007e0000007f000000ff0000007f0";
 when "01111101100" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41500ff800f00ff511700fe000780554007c0000003c011110740000007e0040007400000076011100770000007a0000007c0000007c0010107c000000fe000000fd000000fe000001ff0";
 when "01111101101" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff800e00ff511700fe0007805540074000000780111107c000000fc004000740000006e01110076000000f200000074000000f80010117c000000fc000001fc000000fe000001ff0";
 when "01111101110" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff800e00ff511f00fe000f005540070000000f801111170000000f80040005c000000ec01110174000000f6000001f4000000f8001011f0000001f8000001fc000001fe000001ff0";
 when "01111101111" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff800e00ff511f00fe000f005540070000000f0011111f0000000f800400070000000f80111017c000000f8000001f4000000f0001011f0000001f8000001fc000003fc0000037c0";
 when "01111110000" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff800e00ff511f00fe000f005540070000000f0011111f0000000f0004000f0000000f801110170000000f8000001f0000001f0001011f0000003f8000001fc000003fc0000037c0";
 when "01111110001" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff800e00ff511f00fe000f005540070000000f0011111f0000000f0004000f0000000f001110170000001f0000001f0000001f0001001f0000003f8000001fc000003fc0000037c0";
 when "01111110010" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff801e00ff511f00fe000f005540070000000f0011111f0000001f0004001f0000001f001110170000002f8000001f0000001f0001001f0000003f8000001fc000003fc0000037c0";
 when "01111110011" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff801e00ff511f00fe000e005540070000000f0011111f0000001f0004005f000000ef8011101f0000000f8000001f0000001f0001001f0000003f8000001fc000003fc0000037c0";
 when "01111110100" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41c00ff801e00ff511f00fe000e0055401f0000001f0011113f000001ff0004015d0000000f8011111f0000000f8000001f0000001f0001001f0000003f8000001fc000003fc0000037c0";
 when "01111110101" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41c00ff801e00ff511c00fe001e0055401f0000003e0011157f0000003f0004001f0000000f8011101f0000001f8000001f0000001f0001001f0000003f8000001fc000003fc0000037c0";
 when "01111110110" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41c00ff803c00ff511c00fe001e0055545e00000ffe0011115f0000001f0004001f0000000f8011101f0000001f8000001f0000001f0001001f0000003f8000001fc000003fc0000077c0";
 when "01111110111" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011015f0000001f0004001f0000000f8011101f0000001f8000001f0000001f0001001f0000003f8000001fc000003fc000007fc0";
 when "01111111000" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe02000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011115f0000003f0004001f0000000f8011101f0000001f8000001f0000001f0001001f0000003f8000001fc000003f8000007fc0";
 when "01111111001" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe02000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011115f0000003f0004001d0000000e8011101d0000001f8000001f0000001f0001001f0000003f8000001fc000003f8000007fc0";
 when "01111111010" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011115f0000003f0004001f0000000f8011101d0000001f8000001f0000001f0001001f0000003f8000001fc000003f8000007fc0";
 when "01111111011" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055555c000003fe0011115f0000003f0004001f0000000f8011101d0000001f8000001f0000001f0001001f0000003f8000003f8000003f8000007fc0";
 when "01111111100" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe201e0055555c000003fe0011115f0000003f0004001f0000000f0011101f0000001f8000001f0000001f0001001f0000003f8000003f8000003f8000007fc0";
 when "01111111101" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe201e0055555c000003fe0011115f0000003f0004001f0000000f0011101f0000001f8000001f0000001f0001001f0000003f8000007f8000003f8000007fc0";
 when "01111111110" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe201e0055555c000003fe0011115f0000003f0004001f0000000f0011101f0000001f8000001f0000001f0001001f0000003f0000007f8000003f8000007fc0";
 when "01111111111" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe201e0055555c000003fe0011115f0000003f0004001f0000000f0011101f0000001f8000001f0000001f0001001f0000003f0000007f8000003f8000007fc0";
 when "10000000000" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055555c000003fe0011115f0000003f0004001f0000000f0011101f0000001f8000001f0000001f0001001f0000003f0000007f8000003f8000007fc0";
 when "10000000001" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f8001001f0000003f0000007f8000003f8000007fc0";
 when "10000000010" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055545c000003fe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f8001001f0000003f0000007f8000003f8000007fc0";
 when "10000000011" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511400fe001e0055545c00000bfe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f0000007f8000003f8000007fc0";
 when "10000000100" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511400fe001e0055545c00000bfe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f0000003f8000003f8000007fc0";
 when "10000000101" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe02000ffc41400ff803c00ff511c00fe001e0055545e00000ffe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f8000003f8000003f8000007fc0";
 when "10000000110" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41400ff803c00ff511c00fe001e0055545e00000ffe0011015f0000003f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f8000001f8000003f8000007fc0";
 when "10000000111" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41400ff803c00ff511c00fe001e0055545f00000ffe0011115f0000003f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f8000001fc000003f80000077c0";
 when "10000001000" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41400ff803c00ff511c00fe001e0055405f00000ffe0011115f0000001f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f8000001fc000003f80000077c0";
 when "10000001001" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc41400ff803c00ff511c00fe001e0055405f00000afe0011155f0000001f0004001f0000000f0011101f0000001f0000001f0000001f0001011f0000003f8000001fc000003f80000077c0";
 when "10000001010" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc45400ff803c00ff511c00fe001e0055401f0000007e0011157f0000001f0004001f0000000f0011101f0000000f0000001f0000001f0001011f0000003f8000001fc000003fc000007fc0";
 when "10000001011" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc45400ff803c00ff511700fe001e005540170000003e0011057f000000bf0004001f0000000f001110170000000f0000001f0000001f0001011f0000003f8000001fc000003fc000007fc0";
 when "10000001100" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc45400ff803e00ff511f00fe000f005540070000001f0011157f000003ff0004040f0000000f001110170000000f0000001f0000000f0001011f0000001f8000001fc000003fc000003fc0";
 when "10000001101" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41400ff801e00ff511f00fe000f005540070000000f0011111f000003bf000405470000000f801111070000000f0000001f0000000f8001011f0000001f8000001fc000003fc000003fc0";
 when "10000001110" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc41500ff800f00ff511700fe0007005540070000000f8011111f0000003f80040057800000078011100700000007800000070000000f8001001fc000001f8000001fc000003fc0000017c0";
 when "10000001111" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40540ff800380ff5117c0fe0003805540050000000380111107d000000fc004001fc0000003c0111007c000000380000007c0000007c0010007c000000fe000001fc000001fe000001ff0";
 when "10000010000" => data <= 768x"ffe00000ffd40000ffe000007fd10000ffe00000ffc40150ff8001e0ff5111e0fe0003e0554001c0000003c011110340000003e0040007c0000003e0111001c0000003e0000007e0000003e00100077000000ff000001ff000001ff000001ff0";
 when "10000010001" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffc40050ff8000f0ff5111f0fe0003e0554001c0000003e011110370000003f0040007f0000003e0111001f0000003f0000001f0000003f8010007f0000007f8000007fc00000ffc00001ffc";
 when "10000010010" => data <= 768x"ffe00000ffd40000ffe000007fd10100ffe00000ffd40050ff8000f8ff511170fe0001f0554001c0000001e011111171000003f0040001f0000003f011101170000001f0000001f0000001f8010101fd000003fe000005fd000007ff000007f7";
 when "10000010011" => data <= 768x"fff00000fff40000ffe000007f710100ffe00000ffd40014ffc0003cff51107cff0000f855400070000000f811110171000001f8040001fc000000f8111001f0000000f80000007c000000fe01010177000000ff000001ff000001ff00000177";
 when "10000010100" => data <= 768x"fff00000fff40000fff800007f710100fff00000ffd40005ffe0000eff51101fff80003e5540007c0800003c1111007c0000007e0400007f0000007e1110105c0000003e0000005f0000003f0101003f0000003f0000007f000000ff0000007f";
 when "10000010101" => data <= 768x"fff80000fff40000fff800007f750100fff80000fff40001ffe00003ffd11007ffa0000f5540000f0800000f1111011f0000001f0400001f0000000f111010170000001f000000170000000f0101001f0000001f0000001f0000003f00000017";
 when "10000010110" => data <= 768x"fffe0000fffd4000fffe00007f7d0100fffe0000fffd0000fff8000077f510013fe00001555400010000000115110101000000030400000100000003111000010000000300000001000000010101000100000003000000070000000700000007";
 when "10000010111" => data <= 768x"ffff80007fff4000ffff80007f7f5100ffff80007fff40003ffe00005ffd10002ffa0000555400000080000011110100000000000400000000000000111000000000000000000000000000000101000000000000000000000000000000000001";
 when "10000011000" => data <= 768x"3fffe0005ffff0003fffe0005f7f71003fffe0005fffd0000fffc0001777500003ff0000555540000000000011110100000000000404000000000000111110000000000000000000000000000101000000000000000000000000000000000000";
 when "10000011001" => data <= 768x"0ffff80057fffc000ffff800177f750007fff80057fff4000bfff80015ffd11000ffa000455550000008000011110100000000000404000000000000111110000000000000000000000000000101000000000000000000000000000000000000";
 when "10000011010" => data <= 768x"03ffff0055ffff4003ffff0015ff7f0103fffe00457ffd0000fffe001177f510003ff000445554000000800011111101000000000404000000000000111110000000000000000000000000000101010000000000000000000000000000000000";
 when "10000011011" => data <= 768x"007fffe0557fffd000ffffe0117f7fd1003fff80055fff40003fff801157ff100007fe00045555000000800011111101000000000404040000000000111111100000000000000000000000000101010000000000000000000000000000000000";
 when "10000011100" => data <= 768x"003ffff8045ffff4000ffff8111f7f75000ffff00457fff4000fffe01115f7d10003ff80004555400000080001111511000000000004040000000000111111100000000000000000000000000101010000000000000000000000000000000000";
 when "10000011101" => data <= 768x"0003fffe0055fffd0003fffe01177f7d0003fffe0005fffd0000fff8111177f500003fe0000555540000000001111511000000000004040080000000001111118000000000000000800000000101010180000000000000008000000000000000";
 when "10000011110" => data <= 768x"0000ffff00057fff0000ffff01117f7f0000ffff00057fff00003ffec1115ffde0002ffac0005554e000008071111111f0000000f0000404f000000070111111f0000000f0000000f000000070010101f0000000f0000000f0000000f0000000";
 when "10000011111" => data <= 768x"00003fff00005fff00003fff01115f7f00003fff00045fff00000fff141117773c0003ff1c0015551c0000081d0111111e0000001c0004041e0000001f1111111e0000001f0000003e0000001f0101011f0000001f0000001e0000001f000000";
 when "10000100000" => data <= 768x"00000fff000057ff00000fff0001177f000007ff000015ff000003ff071111ff038000ff07c005550380000801c1111503c0000005c0040403c0000001c0111103e0000001c0000003e000000341010103e0000005c0000003e0000007f00000";
 when "10000100001" => data <= 768x"000003ff000005ff000003ff000115ff000003ff000005ff000000ff0071117700f0003f00700055003800000171111100380000007c000400780000007c111100380000007c0000007c0000007c0101003c0000007c0000007c000000740000";
 when "10000100010" => data <= 768x"000000ff0000057f000000ff0001117f0000003f0000055f0000003f00141117001e000f001f0055000e000000070111000f0000000f0004000f000000070111000f800000070000000f800000170101000f8000000f0000000f800000170000";
 when "10000100011" => data <= 768x"0000003f0000017f0000007f0001117f0000003f0000045f0000003f00071117000f0003000700550003800000070111000380000007c004000780000007d111000380000007c0000007c000000741010007c0000007c0000007c0000007c000";
 when "10000100100" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000001f00071117000780030007c055000380000001c1110003c0000007c0040003c0000001c1110003c0000007c0000003c000000741010003e0000007c0000003e00000075000";
 when "10000100101" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030007c0550001c0000001c1110003c0000001c0040003e0000001c0110003e0000001c0000003e000000341010003e0000001c0000003e0000003f000";
 when "10000100110" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030007c0550001c000000141110003e0000001c0040003e0000001d0110003e0000001c0000003e000000141010003e0000001c0000003e0000001f000";
 when "10000100111" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030005c0550001c000000141110003e0000001c0040001e0000001d0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101000" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030005c0550001c000000141110003e0000001c0040001e0000001d0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101001" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030005c0550001c000000141110003e0000001c0040001e0000001d0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101010" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030005c0550001c000000141110003e0000001c0040001e0000001d0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101011" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f00011117000380030005c0550001c000000141110003e0000001c0040001e0000001d0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101100" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f000151170003c0030005c0550001c000000141110003e0000001c0040001e0000001f0110003e0000001c0000003e000000161010003e0000001c0000003e0000001f000";
 when "10000101101" => data <= 768x"0000003f0000007f0000003f0001117f0000003f0000045f0000000f000151170003c0030005c0550001c000000141110003e0000001c0040001e0000001f1110003e0000001e0000003e000000171010003e0000001e0000003e0000001f000";
 when "10000101110" => data <= 768x"0000003f0000005f0000003f0001115f0000003f0000045f0000000f000151170003c0030005c0150001e000000141110003e0000001c0040003e0000001f0110003e0000001e0000003e000000171010003e0000001f0000003e0000001f000";
 when "10000101111" => data <= 768x"0000003f0000005f0000001f0001111f0000000f00000457000080070001d1150003e0020001c0050001e000000141110003e0000001c0040003e0000001f0110001e0000001f0000003e000000371010003e0000001f0000003e0000001f000";
 when "10000110000" => data <= 768x"0000000f000000570000000f000101170000000300000005000080010003c1110003e0000001c0040001e000000171110003e0000001f0040003e0000001f0110001e0000001f0000003e000000371010003e0000001f0000003e0000001f000";
 when "10000110001" => data <= 768x"000000070000005700000003000101150000000300000005000180000003c1110003e0000001c0040000e0000001f1110003e0000001f0000003e0000001f0110003f0000001f0000001f000000170010003f0000001f0000003e0000001f000";
 when "10000110010" => data <= 768x"0000000300000045000000000001011100000000000140050003c0000003c1110003e0000001f0000000e0000001f1110001e0000001f0000003f0000001f0110003f0000001f0000001f000000170010003f0000007f0000003f0000001f000";
 when "10000110011" => data <= 768x"0000000000000045000000000001011100000000000140050003e000000771110003e0000001f0000000e0000001f1110001f0000001f0000003f0000001f0110003f0000001f0000001f000000170010003f0000007f0000003f0000001f000";
 when "10000110100" => data <= 768x"00000000000000450000000000000111000000000001c0050003e000000771110003f0000001f0000000f0000001f1010001f0000001f0000003f0000003f0110003f0000001f0000003f800000170010003f8000005f0000003f8000007f000";
 when "10000110101" => data <= 768x"00000000000000050000000000000111000000000001d0040003e0000003f1110003f0000001f0000000f000000171010001f0000001f0000003f8000003f0000003f8000001f0000003f8000001f0010003f8000001f0000003f8000007f000";
 when "10000110110" => data <= 768x"00000000000000040000000000000111000020000001f0040003f0000003f1110003f8000001f0000000f800000171010001f8000001f0000003f8000003f0000003f8000001fc000003f8000001f1000003f8000001fc000003f8000007f000";
 when "10000110111" => data <= 768x"000000000000000400000000000001110000e0000001f0040003f800000370110001f8000001fc000000f800000171010001f8000001fc000003f8000003fc000003f8000007fc000003f80000017c000003f8000001fc000003f8000003fc00";
 when "10000111000" => data <= 768x"000000000000000400000000000011110001f0000001f0040003f8000003fc110003f8000001fc000000f80000017d010001f8000001fc000003fc000003fc000003fc000007fc000003fc0000037c000003fc000001fc000003fc000003fc00";
 when "10000111001" => data <= 768x"000000000000000000000000000051110001f0000001fc000003fc000003fc110003fc000001fc000000fc0000007d010001fc000001fc000003fc000003fc000003fc000007fc000003fc0000077c000003fc000001fc000003fc000003f400";
 when "10000111010" => data <= 768x"000000000000000000000000000151110003f8000005fc000003fc000003fc110003fc000001fc000000fc0000007c010000fc000001fc000003fc000003fc000003fe000007fc000007fe0000077c000003fe000001fc000003fe000003f400";
 when "10000111011" => data <= 768x"000000000000000000000000000151010003f8000007fc000003fc000007f4000003fe000001fc000000fc0000007c010000fe000001fc000003fc000003f4000003fe000007fc000007fe0000077c000003fe000001fc000003fe000003f400";
 when "10000111100" => data <= 768x"000000000000000000000000000151010003f8000007fc000003fc000007f4000003fe000001fc000000fc0000007c010000fe000001fc000001fc000001f4000003fe000007fc000007fe0000077c000003fe000001fc000003fe000001f400";
 when "10000111101" => data <= 768x"000000000000000000000000000151010003f8000007fc000007fc000007f4000003fe000001fc000000fc0000017c000000fe000001fc000001fc000001f4000003fe000007fc000003fe0000077c000003fe000001fc000003fe000001f400";
 when "10000111110" => data <= 768x"000000000000000000000000000151010003f8000007fc000007fc000007fc000003fc000001fc000000fc0000017c000000fc000001fc000001fc000001fc000003fe000007fc000003fe0000077c000003fe000001fc000003fe000001ff00";
 when "10000111111" => data <= 768x"000000000000000000000000000150010003f0000007f4000007f8000007fc000003fc000001fc000001fc000001fc000001fc000001fc000003fc000003fc000003fc000007fc000003fc0000077c000003fe000001fc000003fe000003ff00";
 when "10001000000" => data <= 768x"000000000000000000000000000140010003e0000007f000000ff8000017f000000ff8000007fc000003f800000178000001f8000001fc000003f8000007fc000003f8000007fc000007f80000077c000003fc000007fc000007fe000007ff00";
 when "10001000001" => data <= 768x"000000000000000000000000000001010003e0000007f000000ff8000017f000000ff8000007fc000007f8000007f8010003f8000007f8000003f8000007f0000007f8000007f800000ff80000177c00000ffe00001fff00000fff800017ffc0";
 when "10001000010" => data <= 768x"0000000000000000000000000001010100000000000150000003f80000077c110007fe000007fe00000ffe0000077f010003fe000005fc000007fc000007f400000ffc00001ffd00001fff0000177f00003fffe0007ffff000effff801d7f5fc";
 when "10001000011" => data <= 768x"0000000000000004000000000000151100003f000001ffc40001ffc0000177c10003ffe00003ffc00003ffc000077fc10007ff80001fff00003fff00007ff70001ffff8001fffdc007ffffe0077fff703ffffff87dfffffcfbfffffe777f777f";
 when "10001000100" => data <= 768x"0000000000000045000038000001ff110003ff000007ff04000fff00001ff711001fff00001fff00003fff00001ff701003fff00017ffc000ffffe007577fd00c3bfffa0157fffc0383fffe0757f7f70fffffff85ffffffceffffffc77fffffc";
 when "10001000101" => data <= 768x"000000000000005500000000000101110007e000001ff005003ff000007ff11100fff00000fffc0000fff80001777d0100fff80001fff40000fff00001fff00001fff00055fffd00ffffff0077ff7f00ffffff80ddffffc008ffffc001ffffd0";
 when "10001000110" => data <= 768x"00000000000004550000000000011111000000000014004500ff00000177111103ff800007ff400407ff8000077fc1110fffc00007ffc0000fffe00007ffc0000fff80000fff80000fff8000077ff0000ffff80007fffc000ffffe0007ffff00";
 when "10001000111" => data <= 768x"00000002000004550000000000011115000000000000044500000000015011110ff800001ffc00443ffc00007f7c01117ffe00007ffc0004fffe000077f70011fffe0000fffc0000fffc00007f7c0001fffe0000ffffc000ffffe000f7f7f000";
 when "10001001000" => data <= 768x"0000000200000555000000000001111500000002000004550000000000001111000000005d000044ff800000ffc10111ffc00000ffc00004ffc000007ff00011ffe00000fff00000fff000007f700001ffc00000ffc00000ffc00000fff40000";
 when "10001001001" => data <= 768x"000000020000455500000000000111150000000200000555000000000000111100000000000000550000000050010111f8000000fc000004fc000000fc000011fc000000fc000000fe0000007f000001fe000000ff000000fe000fc0fc007ff0";
 when "10001001010" => data <= 768x"000000220000455500000000000111550000000200000555000000000000111500000000000000550000000000010111000000000000000480000000c0000011c0000000c0000500c0001f80c1007fc1e000ffe0c001ffc0e001ffe0c00177f0";
 when "10001001011" => data <= 768x"00000022000055550000000a000111550000000200000555000000000001115500000000000000550000000000010111000000000000000500000000000010110000fe000001ff000003ff0000077f010007ff000007ff00000fff80001fff00";
 when "10001001100" => data <= 768x"00000022000055550000000a00011155000000220000055500000000000111550000000000000455000000000001011100000000000170050001fc00000777110007fe000007fd00000ffe00011f7c01003ffe00007ffc00007ffe00007ffc00";
 when "10001001101" => data <= 768x"0000002b000055550000000a000111550000c8220000dd550000d808000157550000f6020007fd550003fb000001fd150001f8000001f0050003f0000017f111000fe000001fc000003fe000007f710100fff00001fff00001fff000017ff000";
 when "10001001110" => data <= 768x"0000022b00005555000000aa000115550000022a000155550001200a00017155000168220005d5550007e000000775150003f0000007c4550007e0000007c111003f8000007f0000007f8000007fc10101ffe00001ffc00003ffe00007fff000";
 when "10001001111" => data <= 768x"000002bb00055555000000af001115550000022b00055555000000aa00055555000d802200055555000f6000001f5555001fa002001fd555001f8000001f1111001f0000005f004400fe000001fc011103fe000007ff000007ff800017ff0000";
 when "10001010000" => data <= 768x"000023ff0005555f00000aff01115557000003bf0005555500000aaf011155550020023b00445555006800aa00511555007a00220174455500ff000001fd115500f8000001f4445500f8000005f111110fe000001ff000041ff8000017fc0111";
 when "10001010001" => data <= 768x"0002bfff00555fff0000ffff01155f7f00023fff000557ff00002fff011157ff00003bff004555ff00000aff0351557702c003bf07d5555503a000af074115550ff800221fd055550fc0000007c111150f8000001f0004457f00000077001111";
 when "10001010010" => data <= 768x"003fffff055fffff00bfffff115f7f7f003fffff0557ffff002fffff1157ffff002fffff0055ffff000bffff01157f7f0003ffff10557fff2602ffff351557ff29803fff7d0555ff7e800aff7f515557fe00023b7c045555f8000008f0111155";
 when "10001010011" => data <= 768x"3fffffff5fffffff0fffffff577f7f7f2fffffff57ffffff0fffffff57ffffff2fffffff57ffffff0fffffff177f7f7f03ffffff55ffffff02ffffff157fffff22ffffff555fffff68bfffff55577f7fb02fffff5555fffff80affffd1157fff";
 when "10001010100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffff77ffffffffffffff7fffffff3fffffff5f7f7f7f3fffffff5fffffff8fffffff57ffffff";
 when "10001010101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001010110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001010111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffc7fdff3fe7f8ff1f47fc7";
 when "10001100000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffffffffffffe7ffff17c7f5ff1fe7f8ff1fc7fdff9fe3f8ff1fc7f07";
 when "10001100001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffffffffffffeffff717c7f5ff1fe7f8ff1fc7fdff9fe3f8ff1fc7f17";
 when "10001100010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7ffff9fe3fcf71f77fc5f9fe3f8ffdfd1fc7f8fe3f80d1ff3745";
 when "10001100011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fdffcfe3f8f79ff1fc7f8fe0f80d5ff1fc5f8ff3fc7f9f717c7";
 when "10001100100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fdffcfe3f8f79ff1fc7f8fe0f80d5ff1fc7e0ff3fc771f717c7";
 when "10001100101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fdffcfe3fcf71ff1fc7f8fe0f80fdff1fc5e8ff3fc751f737c7";
 when "10001100110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fddf9fe3f8f71ff7fc7f9fe0fc2fdff1fc5f9ff3fc751f737c7";
 when "10001100111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fddfbfe3fcf717f7fc7f9fe1f80fdff07c5f9fe3fc771f777c7";
 when "10001101000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffbffffdff1fcff9ff3fcf717f3fd5f9fe1f82f1ff47c7f1fe3fe711ff3fc7";
 when "10001101001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff7fd7fbff3f8ff1ff1fc7f9fe3fc271ff1fc1f9ff0fc771ff5fc709fe3fe711f71fc7";
 when "10001101010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffff7feff5ff7fc7f9fe3fcff1fc7fc5f9fe3fc0717f5f45f1fe7fe701fc7fc700fe3fc7407e17c7";
 when "10001101011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7ffffffffffdff7fdff9fe7fcff1fc7fc7f9fc7fcff9fc7fc5f9feffc0717c7f4701fe3fcf01fc1fc7c0fe1f87f0757707";
 when "10001101100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffffe7ffffdf47fdff8f87fcffdf477c5f9fe7fc3f9fc7fc1b9fcffcc11fc7fc700fc3f8fc07c1fc7f8fc3f87fdfd7f07";
 when "10001101101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7d7f7f7ff8fa3feffcf57fc7fcf87fcf7dfc77c7f8fe7fc055fc7fc500fc7fcf417c7fc7e0783f87f07c7f07f9febf87f5fff757";
 when "10001101110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffffffffffffffff7ffffefe3fff7d757f57fcf83f8ffc7c7fc7fcfe7f03f5ff7f1520fe7f8f04fc7fdf80fc3f8f707c7f07f87e3f87fdffffc7f9febfaffdfd77f7";
 when "10001101111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffdff7fdffcfe3f8f7c7f7fd7fcf83f8ffdfc7c07f8fe7e9f55f77f1f00fe3f9fc07c7f1ff87c3f0f7c7d7f07f9febfaffdff7f7ffcfebfaff47d7f77";
 when "10001110000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffbffdff7f9ff8fe3f8f7c7f7d17fcf83e1ffdfd7d1fa8fe3f3f047f7f1f807e3f1ff47c1f1ff83c3e0f7d7f7f5ff9febf2ffdfd5f7ffefe3feffc757757";
 when "10001110001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffdfffff7f9ffdfe7f9ff8fe3f8f7d7d7c1ffcf83e1f55fd7f1f00fe3f9f40773f1ff07e3e1ffc7c1c1ffc3e3e0f7d7f7f7ffcfebf6ffc7d5f7ffc7e3f2f557d7717";
 when "10001110010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffdf77f5ffcfe3f8ffcff7dd7fcfe3c0ffd7c3d1ff8fd3f9f147f1f1f807e3f1fd0773f1ff83e3e1ffc7f1f1ffcfebfaf7dff5f7ffefe3f6ffc7f5f5ffc3e3e0f557d7757";
 when "10001110011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffbffff57f17dffcff3f8ffc7f1d57feff1c0ffc7f1f1fb87fbf9f047f1f1fc03e1f0ff03c1717fc3f3e0ffc7f5f5ffefeffef7f7f5f5ffe7f3fffdc7f5f5f8e3fbf8f557ffd57";
 when "10001110100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffff7fdffffeff9ffff47f17dffe7f878ffc7f05dffe7f9c0ffc7fdf1f183f9f9f407f1f1fe03e0f0ff4171f17fe3ffe0ffc7f5f5ffe7effaf7f7f5f5ffe3f8f1f5d5fd71f8e3fff8f557fff57";
 when "10001110101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffff7f5ffffe7f9ffff67f17dffe3f878fff7f55dffe3f9e0f5d7f5f1f003f8f9fc15f1f1ff83f0f0ffc1f571ffe3fff0ffc7f5fdffe7f8fafff7f175ffe3faf0f555ff55f8a3fff8fd57ff757";
 when "10001110110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffff7f1fdffe3f9bcfff7f17d7fe3f878fff7fdd45fe3f9e0f547f1fdf003f8f8fd01f071ff81f8f0ffc1f5717fe3f7f8ffc7f5fdfff7f8fafff7f575fbe3fff0f555fff57c2bfffcff57fffd7";
 when "10001110111" => data <= 768x"ffffffffffffffffffffffff7f7fff7fffffbfffff7f1fd7fe7f9fc7f77f17c7fe3f87c7fc7fdf45fc7f9f43157f1fc7803f8f8ff01f0707fc1f8f0fff5f5f57fe7fffafff7f5fffff3f8fafff3f57178e3fff8fd55fff57e0ffffe3f57ff775";
 when "10001111000" => data <= 768x"ffffffffffffffffffffffff7f7f7f77ffffbfefff7f9fc5fe7f9fe7f47f17c5fe7f83e0fc7fdfc79c7f9fe7057f1f47e03f8fc7f41f0fc7fe1f8f87ff5f5fd7fe7fbfbfff7f5f77ff3f8fafd71fd707823fffe3d55fffd5e0fffffc757ff7f7";
 when "10001111001" => data <= 768x"ffffffffffffffffffffffff7f7f7f77ffffbfe7fd7fdfc5fc7f9fe7747f17d1fe7f87e3fc7f97d7887f9fe3417f1f47e03f0fc3fc1f0fc7fe1f9fc3fe7f5fd7fe7f8fbfff7f5f77ff3f8faf551f5757823fffe3d57fffd5f8fffffff57ffff7";
 when "10001111010" => data <= 768x"ffffffffffffffffffffffff7fff7f77ffff9fe7fc7fdfc7fc7f9fe37c7f17c1fe7f8fe3dc7f97f7827f9fe7417f1f47f03f0fc3fc1f1fc7fe1fbfc3f47f5fd7ff7f0fbfff7f5ff7fe3fcf83555ff757e23fffe3d57fffddf87ffffff57ffff7";
 when "10001111011" => data <= 768x"ffffffffffffffffffffffff7fff5f77feff9fe3fc7f1fc7fe7f9fe37c7f17d1fe7f2fe3547f17f7827f1fe7d07f1f47f03f0f83fc1f5fc7fe7fffc7f77f5fd7ff3f1fbfff5f5fd7ee3faf87575ff757e27fffebf57fffd5f87ffffffd7fffff";
 when "10001111100" => data <= 768x"ffffffffffffffffffffffff7fff3f77fcff3fe7fc7f1fc7fefe3fe7fc7f17c1fc7f3fe2547f1fc7807e1fe7d07f1fc7f83f1f83fc5f5fc7fe7fffcff77f5fd7ff3f3faffd5f5fd7ee3fbfc7557fff57e0ffffe2f57ffff5f87ffffffd7ffff7";
 when "10001111101" => data <= 768x"ffffffffffffffffffff3fff7d7d3f7ffcf83fe7fc7c7fc7fefe3fe7fc7f7fc5fcfe7fe0147e7fc5807e3fcfd07f1fc7f83e3f87fc7fdf07fefeffcff7775fd7ff3e3fafdd5d7fc78e3effcf557f7f55e2ffffe3f57ffff7f87ffffffd7ff7ff";
 when "10001111110" => data <= 768x"ffffffffffffffffffffbfff7d753f77fcf83fe7fc7c7fc7fefe3fe7fc7f7fc1f8fe7fc0147c7fc580fc3fcfd17c1fc7f83e3f87fcffdf07fefebfcfff7d5fd7fe3e3fafdd7d7f478e7fffcf557f7fd7e3fffffbf57fffdff8fffffffdffffff";
 when "10001111111" => data <= 768x"ffffffffffff7ffffffe3fff7d757f57f8f83fc7fcfc7fc5fcfe7fcffd777f51b0fe7f8804fc7fdf80fc3f8fd07c7f07f07ebf0ffdffff07fcfebfaff77d777ffe7e3f3fdc7d7f578effff8f557f7f57e3ffffa3f57fffd5f8fffffffdffffff";
 when "10010000000" => data <= 768x"ffffffffffff7ffffffe7ffff17f7f5ff9fa3f8ffdf47fdff9fe7e0f71fc7d0739fe7f1f15fc7f1f00fc7f1fc07c7f17f07e3e0ffdfd7f5ff8feff7ffd7d7f5ffe7e3f7f5c7d7f5f8cffff8f557f7f5fa3ffff8fd5ffffd7f8fffffff5fffff7";
 when "10010000001" => data <= 768x"ffffffffffffffdffffeffbf777c7f1ff3fe7f1ff1f47f17fbe0781ff1f47d1723fefe3f11fc7f7f00f87e3f017c7c1fe07c7e1ff17d7f5ffbfc7efff5fd7f5ff8fa7eff54757c5f18fffe3f557f775f83ffff3fd5ffff7fe1fffffff5ffffff";
 when "10010000010" => data <= 768x"fffffffffffffffffffbffbf77717f17c7f8ff3fc7fdfd5fe7f0f83fe7d1f47fa3f8fe7f57fcfc7f03f8fc7f11707d7f01f8783fc1fdfc7fe3fafebff7f17df7fbf8ffbfd1f5fd5fa1fff83f777f757f0ffffe3f57fffd7f87fffeff57fff7f7";
 when "10010000011" => data <= 768x"fffffffffffffffffff7feff7f73fc7f3fe3fe3f1ff1fc5f3fe3e07f1fd1707f3fb3f8ff1ff1fcff8fe1f8ff0771f07f07e1f07f07f5f07f8ffdf87f1ff5fd778fe1fb7fc7f5fd7fc7e3f87f57d7717f8ffff27f5ffff57f3ffffcff7ffffdff";
 when "10010000100" => data <= 768x"ffffffffffdffdffffcff8ffff47717fff8ff8ffffc7717fff8620ffff0741f7ff27e1ffffc7f1ffffc7f1ff7fc7f1ff7f83e1ff7f47c1ff3fc7e0ff77d7f1f7ffb3f5ff7fd7f5ff7f87fcff7fd7f5ff3f87e0ff5fd7d5ff7fbfa0ff7f7f75f7";
 when "10010000101" => data <= 768x"ffffffffff7ffffffe3fffff7d1fd77ffe3fc3fffc1fc7fffe1fc3ffff1147ffff1803ffff1d07ffff1f07ff771f477ffe1fc3fffc1fc7fffc1f83fffc1f03f7fe9f03fffddf01fffedfc3ff7d5fd77ffe1f93fffd5fd7fffe0f83ffff5711f7";
 when "10010000110" => data <= 768x"fffffffff7ffffffe3ffbfff417f7f7fe03e3ffff07c1fffe07e1fffc17f1fffe08e3ffff1c417fff8e03ffff1711ffff0e03ffff0551fffe07e1ffff07c1ff7e07c1fffc07c1fffecf80fff6570077feef80fffcdfc1fffe8fe9fffd57c57f7";
 when "10010000111" => data <= 768x"fffffffffffdfffffffbffff37d17f7f23e1ffff05c1ffff0fe0ffff07d1ffff02e0bfff14417fff0e00ffff1d01ff7f0c00ffff1d11ffff0ff0ffff07f17ff703e0ffff01c07fff01e0ffff01c07f7f0f807fff5fc07fffcf807fff5fd07fff";
 when "10010001000" => data <= 768x"ffffffffffdffffffe0fffffff077f7ffe02ffff7f05ffff3f07ffff7707f7ff7807ffff1407ffff0807ffff11077f7fc303ffffc707ffffff83ffff77c3ffffff83ffff7f05ffff3f03ffff1f017f7f1e03ffff5c01fffff803fffff001ffff";
 when "10010001001" => data <= 768x"fe1fbffffc1d7ffff80bffff7c17ff7ffc07fffffc01fffff801ffff1001ffff1003ffff1007ffff800fffffc4077f7fbe07ffffff07fffffe07fffff707fffffe07fffffc07fffffc07ffff7c077f7ff803fffff007fffff003ffff7007ffff";
 when "10010001010" => data <= 768x"f80fbffffc0d7ffff80bbfff7c15177ff8001ffff4001fffe0003fff710177ffe003ffffe007ffffe007ffff77077f7fff07ffffff07ffffff07ffffff07f7fffe03fffffe07fffffe03ffff7c037f7ffc03fffffc01fffff801fffff001ffff";
 when "10010001011" => data <= 768x"ff3ffffffc0ffffffc0fafff7517177f80001fffc4011fff8e023fffc5017fffe0007fffc005ffffe007ffff7d077f7fff03ffffff07ffffff03ffffff07ffffff03ffffff07fffffe03ffff7f017f7ffe01fffffc01fffffc00fffffc007fff";
 when "10010001100" => data <= 768x"ff07fffffc07fffffe07ffff7407d77ff00383ffd00447ffe3008ffff10117fff0003ffff0017ffff003ffff77037f7fff83ffffff01ffffff83ffffff077fffff83ffffff01ffffff01ffff7f01ff7ffe01ffffff01fffffe00fffffc007fff";
 when "10010001101" => data <= 768x"ff03ffffff01fffffe03ffff7f017f7fff03bfffff0155fffe0000fff700107ffe00017ffc0005fffc018fff7d01ffffff81ffffffc1ffffff81ffffffc1ffffff81ffffff01ffffff80ffff7f017f7fff00ffffff007fffff007ffff70077ff";
 when "10010001110" => data <= 768x"ffefffffffc5ffffff80ffff7f01ff7fff81ffffffc1f5ffff80effff7c15fffff803fffff40157fff80003f7f00005ffe0080ffff41d7ffffc0ffffffc1f7ffff81ffffffc1ffffffc0ffff7fc17f7fff807fffffc07fffff803fffff001fff";
 when "10010001111" => data <= 768x"fffbfffffffd7ffffff03fff7f517f7fffe03ffffff05dffffe03ffff7f077fffff03fffffd015dfffc0000f7f410507ff80203bff10757fffb03ffffff077f7ffe07ffffff07fffffe07fff7f707f7fffe03fffffc01fffffe03fffffc01fff";
 when "10010010000" => data <= 768x"fffe7ffffffc5ffffff80fff7f701ffffff80ffffffc0d7ffff80bfffff417ffffe0009fffc00107ffc002037fc0011fff80183fffdc1dfffff81ffffff41ffffff83ffffffc1ffffff81fff7f701f7ffff80ffffff007fffff807fffff007ff";
 when "10010010001" => data <= 768x"ffffaffffffc07fffffc07ff7f7d07ff7ffe07ff7dfc055f78e8003f7455007f7c78007f7d50017fff0003ff7f1517ffffbe0ffffffc1ffffffc0ffffffc1ffffffc1fff7ffc1ffffffc0fff7f7c077f7ff803ff7ffc01ff7ff801ff77fc01ff";
 when "10010010010" => data <= 768x"ffff83ffffff01fffffe03ff7f7c017f7ffe03bf5fff017f1ffe03ff375417ff3f1c03ff1f1801ff1f8003ff1743077f3fe607ff7ff707ff3ffe0fff3ff707ff3ffe07ff1fff07ff3ffe03ff1f7c037f1ffe03ff1ffc01ff0ffc00ff1ffc007f";
 when "10010010011" => data <= 768x"fffff1ffffffc07ffffee07f7f7c00753ffe007b1fff005f0fff00ff1ff5017f0fe380ff07f1007f0ff800ff077c417f0ff881ff1ffdc1ff0fff81ff17ffc1ff0fffc1ff07ffc1ff07ff80ff077f017f07ff00ff07ff007f03ff003f01f7007f";
 when "10010010100" => data <= 768x"ffffffbffffffd5ffffffc0fd77f7007efffe00ec7fff00583fff00f03f7701783ff100fc1ff1007c3ff800f01ff001701ff881f01ffd01f01fff83f41fff01fe1fff83fc1fffc1fe0fff81fc1ff711f80fff00fc1fff01f80ffe00f007fc007";
 when "10010010101" => data <= 768x"fffffff3ffffffc1ffffff807d7f7f01f8ffff80f07fff41f83ffe00f07f1501f83f8e00fc7fd400c03fe000401f7101003fff83441fff010c3fff835c1ff701fe3fff83fc1fff01fc1fff01f41f7f01f81ffe01f01fff01f01ffe00f01ffc00";
 when "10010010110" => data <= 768x"fffffffffffffffcfffffff87fc77f70ff83fff8ff07fff0ff83fff8f707f7f0ff83e3b0ff01c140ff01f8807f01fc00ff00fe30ff41fff0ffc3fff8ffc1ff70ffe3fff8ffc1fff0ff81fff0ff017f70ff01ffe0ff01ffc0fe01ffc0fc01ffc0";
 when "10010010111" => data <= 768x"ffffffffffffffffffffffff7f7d777ffff87bfffff051fffff001fff7f057fffff80ffffff0077ffff0063e7f701715fff83f80fffc7fc5fffc3feffffc7ffffff83ffffffc1ffffff83fff7f701f7ffff03ffeffc01ffcffc01ffcffc01ffc";
 when "10010011000" => data <= 768x"ffffffffffffffffffffffff7f7f7fffffffbffffffc1f7ffffc183f7ffc117ffffe01fffffc11fdfffe00f87f7c017dfffe0ff8ffff077cffff0ffcffff07f7ffff0fffffff07fffffe07ff7f7f077ffffe07fffffc07fffffc03fffffc01ff";
 when "10010011001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffbfff7fffc7f7ffff87e77fff0707ffff823f7fffc45fffff803f7f7f001fffff81bfffffc1ffffffe1ffffffc1ffffffe3ffffffc1ffffffc1ff7f7fc1ffffff80ff7fffc1ff7fff80ff7fff0077";
 when "10010011010" => data <= 768x"ffffffff7fffffff7fffffff7f7f77ff1ffff3ff1ffff07f3fffe0ff1ffff0771ffff0ee1ffff1443fffe0061f7f70073ffff0075ffff0573ffff87f7ffff07f3ffff87f7ffff07f3ffff07f1f7f707f1ffff03f1ffff01f0fffe03f07fff017";
 when "10010011011" => data <= 768x"ffffffffffffffffbfffffff1f7f7f7f1fffffff07ffff7f07fffe1f07fffc1f07fffe1f07fffc1f07fffc3f077f7c110ffff80007fffc0107fffe0107fffc1507fffe1f07fffc1f07fffc3f077f7c1f07fffc0f05fffc1f03fff80f01fffc07";
 when "10010011100" => data <= 768x"fffffffff7fffffff3fffffff37f7f7f83ffffff01fffff780ffffc301ffff4180ffff83c0ffffc1c0ffff83517f7f05e1ffff00c1ffff0080ffff8011ffff0080ffff8300ffff0700ffff8f017f7f0700ffff03007fff07007ffe03007fff01";
 when "10010011101" => data <= 768x"fffffffffdfffffffeffffff7c7f7f7fe07ffffbf05ffffde03ffff8f03ffff0f03fffe0f01ffff0f83fffe07c7f7f71f83fffe0f01fffc0e01fffe0f017ffe0e03fffe0001fffc1001fffc3001f7fc1000fffc0001fffc1000fff800007ffc0";
 when "10010011110" => data <= 768x"ffffffffffdfffffff9fffff7f1f7f7df80ffff9fc07fffdfc0ffff0f407fff0fe07fff0fe07fff0fe0ffff87f177f70fe07ffe0fc07fff0fc0fffe0fc07fff1f007ffe14007fff1800fffe000077f600000ffe00001ffc00000ffe00001fff0";
 when "10010011111" => data <= 768x"fffffffffff7ffffffe7ffff7f477f7fff03fffdff01fff4ff83fff0ff01fff0ff81fff8ffc1fff0ffc3fff87f017f70ff83fff0ff01fff0ff03fff0ff01ff71fe03fff05505fff00003ffe001035f7000000fe000001ff080000fe0f0001ff0";
 when "10010100000" => data <= 768x"fffffffffffdfffffff9ffff7f71ff77ffc0fff3ffc07ff0ffe0fff8ffc07ffcffe07ff0fff07ff4fff0ffe07f407f70ffe0fff8ffc07ffcffc0fff8ffc07ff0ff00fff85441fff40001fff80101f771000003f0400001f0e00003f07d0007f0";
 when "10010100001" => data <= 768x"fffffffffffdfffffffeffff7f7c7f7ffff87ffbfff05ff1fff03ff0fff037f4fff03ff8fffc1ffdfffc3ff87f747f70fff03ffefff07ffcffe03ffe77f077feffc03ffe5f107ffc00207ffc00007ffc0000387840000070e8000070fd000070";
 when "10010100010" => data <= 768x"ffffffffffff7ffffffe3fff7f747f7ffff81ffcfff81ffcfff81ff8fff01ffffff81ffefffc1ffcfffe3ffc7f781f7dfff81ffffff01ffffff01fffffd01fffff801fff5d101fff00203ffe01007fff00003ffe0000141ce0000038f4000010";
 when "10010100011" => data <= 768x"ffffffffffff7ffffffe3fff7f7f7f7ffff83ffffff01ffffff81ffffff01ff5fff80ffcfffc1ffcfffc0ffe7f7c1f7ffff81ffefff01ffffff01ffffff01ff7ffe01fffdf141fff08380fff01511f7f00003ffe00001fdc8000020cd000001c";
 when "10010100100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffe3ffffff45ffffff81ffff7f01ffffff81ffffff01ffffff80ffe7f7c1f7dfffe3ffefffc5ffffff81ffffff01ffffff00fffffc01fffbe080fff145c177f00300fff00001fff00001ffe00001554";
 when "10010100101" => data <= 768x"ffffffffffffffffffffffff7f7f1f7fffff8ffffffd1ffffffc07fff7fc07fffffc07fffffc07fffffc07ff7f7d077fffff0ffffffd1ffffffc0ffffff407f7ff3007fffc0007ffffa80fff1ffc077f03f80fff00500fff00000fff00001fff";
 when "10010100110" => data <= 768x"ffffffffffffffffffffefff7f7fc77fffff83ffffff07fffffe03ffffff01ffffff03ffffff01fffffe03ff7f7f037fffff03ffff5f07fffe0c03ffff1403ffffc003ffffc407fffffc07ff1f7c07ff0ffe07ff015c07ff00000fff000017ff";
 when "10010100111" => data <= 768x"fffffffffffff7ffffffe3ff7f7fc17fffff83ffffff01ffffff01ffffff01ffffff03ffffff01fffff201ff7f7701ffffef83ffffc705ffffcc01ffffc001ffffc001ffffd401fffffe03ff5f7c03ff0ffe03ff05fc07ff002807ff000007ff";
 when "10010101000" => data <= 768x"ffffffffffffd7ffffffc3ff7f7fc7ffffff83fffffc01fffffe01fff7ff01ffffff01ffff7f01fffe3f00ff7f1f017fff1f83ffff1f41ffff8c00fff7d0007fff8000ffffc5007ffffe00ff5f7f007f07ff00ff057f00ff002e00ff010001ff";
 when "10010101001" => data <= 768x"fffffffffffff5ffffffe0ff7f7f717fffffe03fffff407fffff007ff7ff0077ffffc03fffffc01fffffc03f7d7fc03ffe0fe07fff07d07fff8f000fffc5001fffe0000fffc0401fffe3c00f7777401f03ffe00f017fc007000fe00f00014017";
 when "10010101010" => data <= 768x"fffffffffffffd5ffffffe0f7f7f7f17fffffe03fffffc01fffff803fffff001fffff803fffffc01fffffc017f777c01ffb3fc03ff407d07ffe0fe03fff07000fff86000fffc0000fffe00007fff1400fffffe00547fff00000ffe0000057f00";
 when "10010101011" => data <= 768x"fffffffffffffff5fffffff87f7f7f75fffffff8fffffff0ffffffe0ffffffc0ffffffc0ffffffd0ffffffe07f7fff70ffffbfe0ffff17f0fff803f8fff503f0ffffe380ffffc100ffffe0007f7ff000fffff030fffff5f0ffeffff8f5037ff0";
 when "10010101100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffff7fffffffffffffeffffffffffffffff7f7f7f7ffffffffffffffdfffffffcfffffff01ffffff80ffffffd1dffffff0c7f7f7f00ffffff80ffffff41ffffffc3fff77ff7";
 when "10010101101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffff7ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffeffffffff5ffffff00ffffff40fffffff87f7f7f70fffffff8fffffffcfffffffcfffffff4";
 when "10010101110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffd017ffff8003ffff0001f4ff8000fe7f00017fff0000ffff0001fffe00003ff000001f";
 when "10010101111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffffffffffffffff7f75577fffe003ffffc001ffff8001ffff00017ff000000ff0000007e000000f70000017f800003ffd00005fff0000ffff000077";
 when "10010110000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7fff7fffffffffffffffffff83fff7f70177ffc00003ffc00001ffc00003ffc000077fe00003fff00017fff8000ff7f0001ffff8000ffff4001ffff8001ffff80017f";
 when "10010110001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7ffffffffffffff45ffffee00ffffc00007ffe00003ffc00007ffe00003f7f00007fff0000ffff0001ffff8000ffff00017f";
 when "10010110010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffff00fffffc007ffff8002fff400001ff800001ffc00001ffc00003f7f00007fff0000ffff0001ffff8000ffff00017f";
 when "10010110011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7ffff00fffffc007fffe0002bff000001ff800001ffc00001ffe00003f7f00007fff0000ffff0001ffff8000ffff00017f";
 when "10010110100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffffffffffffffffffffffffffff7ff017fffff003fffd40015ff800000ff400001ffc00003ffc00001ffe00003f7f00007fff0000ffff0000ffff8000ffff40007f";
 when "10010110101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffaffffff40177fff800fffff0007fff80007f7f00007fff00003fff00007fff80007fff00007fff80003fffc0007fffc0007f7f50007fffe0003fffc0007fffe0007ffff0007f";
 when "10010110110" => data <= 768x"ffffffffffffffffffffffff7f75077fffe001ffffc0007fffe0007fff000077ff80003fff40001fff80003f7f00007fff80003fff00001fff80002ff7f0007fffe0003fffe0007fffe0003f7f70001ffff8003ffffc005ffffe003ff7f4057f";
 when "10010110111" => data <= 768x"ffbfbfffff0405ffff0000ff7f00007fff80003fff40051ffee0031fff40071ffff00f0ffff01f1ffff81f9f7ffc1f47fffe3f87fffe7fc7ffffff9ff7fff7dfffffffbfffffffdfffffff9f7f7f7f9fffffff8fffffffffffffffffffffffff";
 when "10010111000" => data <= 768x"f020000fc0400407e0600207e0400707f0e00303f0400707e0600607f0701707e0f81f03c1fc1f01e0fe3f81f17f7f01f9ffff80fdffff05ffffff8fffffff07ffffff87ffffff07ffffff877f7f7fc7ffffffe3ffffff57ffffff03ffffff17";
 when "10010111001" => data <= 768x"000000000000000000000000004000000020020000600400006006000070040000781e00007c1f0000fe3f00017f7f00a0ffff00c1ffff00c0ffff0001f7ff0080ffff00c1ffff40e3ffffe075ff7f30e8ffff30f47fff10eeffffe0d777f770";
 when "10010111010" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000000070040000780e00007c1f0000fe3f00007f7f0000ffff0001ffff0000ffff0000ffff0000ffff0001ff7f0003ffff8007ffffc008ffff300077ff10";
 when "10010111011" => data <= 768x"000000000000000000000000000000000000000000000000000000000070070000700e0000701f0000f83f00017c7f0000fe7f8001ffff0000ffff8001f7ff0000ffff0001ffff0000ffff8001ff7f0003ffffc005fffff008ffff900077ff10";
 when "10010111100" => data <= 768x"000000000000000000000000000000000000000000000000000002000070070000700e0000701f0000f83f00017c7f0000fe7f8001ffff0000ffff8001f7ff0000ffff8001ffff0000ffff8001ff7f0003ffffc007fffff008fffff0007fff10";
 when "10010111101" => data <= 768x"00000000000000000000000000000100000001000010050000180f80001c1fc0003e3f80007f7fc0007f7fc0007f7fc0007fffc0007fffc000ffff800077ff8001ffff8007ffff000fffff80057f7f5000ffffa0007fff1000ffff000077ff00";
 when "10010111110" => data <= 768x"000003e0000007e000000fe000001fc000007fe00001ffc00003ffe0000777c0001fffc0001fffc003ffffc0017f7fc0003fff80007fff40007fff800077ffc0003fff80001fffc0000fff80001f7f00000fff800007ff000007ff000007f7c0";
 when "10010111111" => data <= 768x"00003fe000007fc00000ffe000017f400007ffc00007ffc0000fffc0015fffc003ffffe0007fffc0003fffc001777fc0003fffc0001fffc0000fffc00007ff50001fff90001fffc0000fffc000077f0000003f00000005000000000e0000001f";
 when "10011000000" => data <= 768x"0003fff00007fff0000ffff0001f7f70001ffff0041ffff007fffff005f7f7f000fffff001fffff000ffffe0017f7f7000ffffe0007ffff0003c3ff0001015f4000000e600000044000000200000001100000000000000000000000300000007";
 when "10011000001" => data <= 768x"00fffffed5fffffcfffffffe7f7f7f7c1ffffffe0ffffffc0ffffffc1ff7f7f41ffffff81ffffffc0ffffffc07ffff7c03aa3bfc010001fc000000ff0000007d0000003800000010000000180000001400000018000001140000008000000145";
 when "10011000010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7f23ffff83001d740000080000010001002bc003f27fc001fd7f8001ff770001ff3f8000ff1f0001ff1f8000ff1f00017f";
 when "10011000011" => data <= 768x"ffffffffffffffffffffffff7fffff7ffffffffffffffffffffffffffff7f7ffffffffffffffffffffffffff7f7f7f7fffffffffd5ffffd7803c3e00001010000000000005c001403fc001f87fc001ffff8000ffff0001ffff8000ff7f00007f";
 when "10011000100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffffffffffffffff7f7f7f7ffffffffffffd5ffffff80fffff100177fe00003ffc00001ff800000f70000017e000000fc1000007e1800007c1100007";
 when "10011000101" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffffffffffffffff7f7f7f7ffffffffffffd5fffffc80bffff0001ffff00007fff00007ffe00003f7c00003ffe00003ffc00001ffc00003ffc00001f";
 when "10011000110" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7fffffffffffff7fdffffe200ff7f40007fff80003fff00001ffe00000ffd000007fe000007fc000007fe0000077d000007ff800007ffc00057ffc0003fffc0007f";
 when "10011000111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffe3ffffffc1ffffff80ffffff001ffffe000ffffc0007dff80007f7f00007fff00003fff00001fff80003fff50001fffe0003fffc0001fffe0003f7f70001ffff0001ffff4001ffffe003fffff001f";
 when "10011001000" => data <= 768x"ffffffffffffffffffe1ffff7f40777fff0003ffff0001ffff8000ffff400077ffc0003fffc0017fffe003ff7ff0077ffff00ffffff01ffffff80ffffff01d7ffffbbe1ffffffc1ffffffc0f7f7f7c07fffffe07ffffff1fffffff0ffffff717";
 when "10011001001" => data <= 768x"ffe03ffffff005ffffe003ff77f0077ff3f007fff1f00fdfe0f80f8ff1701f17e0f81e07c07c1c07e0781c07707c1c07e0383803f51d5c07ffbff803f71ff007ff3ff803ff7ffc07fffffe037f7f7f01fffffe01ffffff05ffffff07fffff707";
 when "10011001010" => data <= 768x"01f003c300f007c100f00f810071170100780f00007c1f0000381e00001c1c0000383800001c1400001c3800401c3000e01e3800f41df000f80ff800f01ff400f03ffc00f07ffc00f87ffe007c7f7f00fc7ffe00fc5fff00f87ffe00f17fff00";
 when "10011001011" => data <= 768x"000000000000000000000000000000000080000001d0000001f0000001f0001000f803a0007c17f000381ff0001c1f70001c3800001c1000001c3800001d7000000ff000001ff000003ff800003f7c00003ffe00007ffc00007ffe000077ff00";
 when "10011001100" => data <= 768x"00000000000000000000000001000000000000000100000003e0000003f0000003f80f00057c1fc000381fe0001c1d70001838f0001c1c70001cb800001ff100001ff800001ffc00003ffc00007f7c00007ffe00007fff00007ffe00007fff00";
 when "10011001101" => data <= 768x"00000000070000000f80000007c0000007e0000007f0015003f003f80170077900781ff8007c1d5000381800001d1d01001c3800001c1800001c3800001ff000001ff800001ffc00003ffc00007f7c00007ffe00007fff00007ffe00007fff00";
 when "10011001110" => data <= 768x"007c0000007c0000007c0000007c0055003e00ff001c05fd001e07f8001607d0001e0e00001c1c00000e1c0000171c00000e180000075c00000ff800001ff400003ffe00007ffc00003ffe00007f7f00003fff00007fff00007fff00007ff700";
 when "10011001111" => data <= 768x"003e0ff0001c1f40000e1e0000171d01000f1e0000071c0000071c0000071c00000338000007fc00000ffc00001ff700003fff00001fff00003fff80007fffc0003fff80001fffc0000fff80001f7fc0001fff800017ffc0001fff800017f780";
 when "10011010000" => data <= 768x"01fb8000007dc000001f80000007c000000780000007d000000ff800001fff00003fff00007fff00007fff80007f7f00003fff80001fffc0000fff80001fffc0000fff800007ffc00007ffc000057fc00007ffc00007ffc0000fffe0001ffff0";
 when "10011010001" => data <= 768x"00ff0000005f0000000f800000070000000380000007f000000ffc00001ff700003ffe00007fff00007fff80007f7f00003fff80001fffc0000fff800017ffc00007ffc00007ffc00003ffc000037f400003ffe00007ffc0000fffe0001ffff0";
 when "10011010010" => data <= 768x"001f80000007c000000380000003c0000003a0000007f400000ffc00001ff500003ffe00005fff00003fff0000177f00000fff000007ff00000fff800007ff000003ff800001ff000003ff8000077f000007ff800007ffc0000fffc0001fffc0";
 when "10011010011" => data <= 768x"000f80000007c000000380000001c0000001c0000005f000000ff800001ffc00001ffe00001ffc00000ffe0000077f000007fe000007ff000003fe000001f7000003fe000001ff000003fe0000077f00000fff00000fff00000fff80001fff00";
 when "10011010100" => data <= 768x"003f8000005dc000000f80000107c100000180000001c0000003f0000007f400000ff8000007fc000007fc0000077c000003fc000001fc000001fc000001fc000003fe000001fc000003fe0000077f000007ff000007ff00000fff00001ff700";
 when "10011010101" => data <= 768x"0003000000110000003980000017c000000380000001c0000001e0000007f0000007f8000007f8000003f800000179000001f8000001fc000001fc000001fd000003fc000007fc000007fe0000177e00001ffe00001dfc00003bfe000011fc00";
 when "10011010110" => data <= 768x"0000000000040000000e00000007010000070000000500000001c000000370000003f0000005f0000003f000000170000001f0000051f0000033f8000037f000003ff800001dfc000003fc0000017c000003fe000001fc000003fe000003fc00";
 when "10011010111" => data <= 768x"00000000000000000000000000010000000180000000500000005000000170000001f0000001f0000007f0000007f0000003f0000005f0000003f0000003f0000003f8000001f0000001f80000017c000003fc000001fc000001fe000001fc00";
 when "10011011000" => data <= 768x"0000000000000000000000000000000000002e0000005c0000006000000070000000f0000001f0000001f8000001fc000001f8000001f0000003e0000007f000000fe000000dc0000009e000000570000003f8000001f0000001f8000001d000";
 when "10011011001" => data <= 768x"00000000000000000000000000000000000020000000500000004000000050000000f2000000f7000000f300000077000000f8000001f4000001f8000001f1000001f0000001f0000003f8000003fc000003f800000170000000380000007000";
 when "10011011010" => data <= 768x"000000000000000000000000000000000000000000004400000028000000140000003e0000001c0000003c0000001c0000003c0000007c0000007e000000750000007e0000007c000000fe0000007c0000001c0000001c0000001c0000001400";
 when "10011011011" => data <= 768x"00000000000000000000000000000000000000000000110000000a000000140000002f000000470000006f0000007f0000000f000000070000000780000017c000000780000007c000000f8000001740000007000000050000000d0000001500";
 when "10011011100" => data <= 768x"000000000000000000000000000000000000000000000500000007000000010000000380000001c0000183c000017740000003c0000001c0000003e0000001e0000003e0000001f0000003e000000750000003c000000740000006c000000440";
 when "10011011101" => data <= 768x"0000000000000000000000000000000000000000000005000000038000000140000001e0000001c0000000e000017770000003e0000001f0000000f0000001f0000001f0000001f0000003f800000170000001a0000001400000032000000340";
 when "10011011110" => data <= 768x"0000000000000000000000000000000000000000000001400000038000000140000000e0000001f0000000e000007770000003f000000070000000f800000170000000f8000001f0000001f800000170000001b0000001300000012000000130";
 when "10011011111" => data <= 768x"0000000000000000000000000000000000000000000001400000008000000040000000e000000070000000f000007770000002f0000000700000007800000070000000f8000000fc000000f800000170000000b0000001d0000001b000000110";
when others => data <= 768x"0";
end case;
end if;
end process;
end;
