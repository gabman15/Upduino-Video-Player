library IEEE;
use IEEE.std_logic_1164.all;
entity rom is
port(
clk : in std_logic;
addr : in std_logic_vector (7 downto 0);
data : out std_logic_vector (767 downto 0)
);
end rom;
architecture synth of rom is
begin
process(clk) is
begin
if rising_edge(clk) then
case addr is
 when "00000000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000100" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00000111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001000" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001001" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001010" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001011" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001100" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001101" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001110" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00001111" => data <= 768x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
 when "00010000" => data <= 768x"000000010000000100000000000000010000000100000001000000010000000100000001000000010000000100000001000000030000000100000003000000030000000300000001000000000000000000000000000000000000000000000000";
 when "00010001" => data <= 768x"0000000000000000000000000000000000000000000000000000000000000000000000080000000c00000008000000050000000f000000170000001f0000001f0000000f00000007000000030000000300000003000000010000000100000001";
 when "00010010" => data <= 768x"0000003f0000005f0000003f0000001f0000003f0000001f0000001f0000001f0000003f0000001f0000003f0000007f0000003f0000005f0000003f0000007f0000003f0000005f0000003f0000001f0000003f0000001f0000000f00000017";
 when "00010011" => data <= 768x"00000fff00000fff00000fff000007ff00000fff00000fff00000fff000017ff00000fff000007ff00000fff0000077f00000fff000007ff000007ff000001ff000001ff000000ff000000ff0000007f0000007f0000007f0000003f0000001f";
 when "00010100" => data <= 768x"000003ff000005ff000003ff0000077f00000fff00001fff00001fff000015ff000003ff000001ff000003ff0000017f0000007f0000001f0000001f0000001f0000001f0000001f0000000f0000001f0000000f000000070000000300000011";
 when "00010101" => data <= 768x"000000ff000001ff000001ff0000017f000003ff000007ff000003ff4000007f400000ffc000007f8000003f0000001f0000000f0000000700000007000000070000000700000007000000070000000700000003000000010000000000000000";
 when "00010110" => data <= 768x"f000007ff000007ff000007ff000007fe000007ff000007fe00000fff010017fe020007fd000007fe000003fc000001fe000000fc0000007c0000007c00000078000000700000007000000070000000700000003000000000000000000000000";
 when "00010111" => data <= 768x"f800000ffc00005ffe00003fff00003ffe00003ffc40007ffe00003ff400007ffe00003ffc04007ffe00007ffc00007ffe00003ffc00001ff800000ff0000007f0000007f0000007e0000007c0000007c0000003c00000008000000010000000";
 when "00011000" => data <= 768x"ff00000fff00001fff80003f7f00001fff80003fff00001fff80003fff100017ff80003fff00001fff80003f7f00001fff80000fff000007ff000007ff000007fe000007fc000007f800000370000001f8000000f0000000e0000000f0000001";
 when "00011001" => data <= 768x"ff80001fffc0001fffe0003f7f40001fffc0003fffc4001fffc8003fffc0001fffc8003fffd0005fffc0000f7fc00007ffc00007ffc00007ffc00007ffc00007ff000003ff000005fe0000007f000000fe000000fc000001fc000000fc000000";
 when "00011010" => data <= 768x"fff0001ffff0001ffff0003f7f70001fffe0003ffff0007fffe0003fff700017ffe0003ffff4001ffff0000f7f700007ffe00003fff00007ffe00003ffc00007ff800003ffc00000ff8000007f000001ff800020ff000040ff000020ff000040";
 when "00011011" => data <= 768x"fff0000ffff00007fff8001f7f70001ffff8003ffffc001ffff8003ffff00077fff8003ffff0001ffff8001f7f700017fff80007fff00007fff00007ffd00007ffc00007ffc00005ffe000017f400001ffc00003ffc00001ff800003ff000041";
 when "00011100" => data <= 768x"ffe0003ffff0001ffff8003f7f71007ffff8003ffffc007ffffc003ffff4003ffffc003ffffc007ffff8007fff71001ffff0001ffff0001fffe0001fffc0001fffc0000fffc00007ffe000077fc00007ff80000fffc00007ff800007ff000007";
 when "00011101" => data <= 768x"fff000fffff0007fffe000ff7f7001fffff800fffffc007ffff8007ffff4007ffff800fffff0007fffe000ffffc0007fffe0007fffc0007fff80007fff000017ff80001fffc0041fff80063f7f00041fff80061fff00041ffe00060fff000417";
 when "00011110" => data <= 768x"ffe000ffffc001ffffc001ff7f70017ffff003fffff001fffff801fffff001f7fff001ffffd001ffffc001ff7fc001ffff8000ffffc0007fff80007fff00007fff80007fff00107fff00083f7f00117ffe00083ffe00107ffe00083ff4001017";
 when "00011111" => data <= 768x"ffa000ffffc001ffffc003ff7fc0037fffe003fffff007ffffe007fffff007fffff003fffff007ffffc003ffffc001ffff8001ffffc001ffff8000fff700007fff00007fff00007ffe00007f7f00117ffe00007ffc00107ffc00007ff000107f";
 when "00100000" => data <= 768x"ff8001ffffc001ffffe003ff7fc0077fffc007ffffc007ffffe00fffff5007ffffe00ffffff007ffffe00fffffc007ffff8003ffffc001ffff8001fff70001f7ff0001ffff0005fffe0000fffc00007ffc0020fffc00007ff80000fff000007f";
 when "00100001" => data <= 768x"ff8003ffffc007ffffc007ff7fc0077fffe00fffffc01fffffc00fffffc01fffffe01fffffc01fffffc00fff7f0017ffff800fffff0007fffe0003fff70003f7fe0003fffc0001fffe0001fffc00017ffc0001fffc0001fff80000fff0000177";
 when "00100010" => data <= 768x"ff0007ffff4007ffff800fff7f001f7fff801fffffc01fffffc01fffffc01fffffe03fffffc01fffff801fff7f001f7fff800fffff0007fffe000ffff70007f7fe2003fffc4007fffe2003ff7c00037ff80003fff84001fff80003fff00001ff";
 when "00100011" => data <= 768x"ff000fffff401fffff800fff7f001f7fff803fffffc07fffffc03fffff4037ffffc03fffffc03fffff803fff7f001f7fff001fffff001ffffe000ffff70017f7fe200ffffc4007fffe2007ff7c00077ff80003fffc4007fff80003fff00001f7";
 when "00100100" => data <= 768x"ff000fffff001fffff801fff7f001f7fff803fffffc07fffffc07fffffc077ffffc03fffffc07fffff803fff7f003f7fff803fffff001ffffe000ffff7001ff7ff000fffff0007fffe0007ff7c00077ffc0003fffc0007fff80003fffc0003f7";
 when "00100101" => data <= 768x"ff800fffff0007ffff800fff7f401f7fffc03fffffc01fffffc03fffffc07fffffc07fffffc07fffffc01fff7fc01f7fff800fffff000fffff800fffff1007f7ff800fffff1007ffff0007ff7f10077ffe0003fffc0007fffe0003fffc0003f7";
 when "00100110" => data <= 768x"ff8007ffffc007ffffc00fff7f701f7fffe01fffffc01fffffe03fffff407fffffe03fffffc01fffffc00fff7f40177fff800fffffc007ffff880fffffc007f7ff8807ffffc407ffff8803ff7f00017fff0003ffff1001ffff0003ffff1001ff";
 when "00100111" => data <= 768x"ffc007ffffc007ffffe00fff7f701f7ffff00ffffff01ffffff01ffffff01fffffe03ffffff01fffffe00fff7fc0077fffc007ffffc007ffff8007ffff9007f7ff8003ffffc401ffff8001ff7fc401ffff8001ffffc401ffff8001ffffd001ff";
 when "00101000" => data <= 768x"fffb07ffffc007ffffe007ff7f70177ffff00ffffff007fffff80ffffff01ffffff01ffffff01ffffff00fff7f70077fffe007ffffc007ffffc003ffffd003f7ffb003ffffd001ffff8000ff7f40017fffa000ffffc001ffffe000ffffc001ff";
 when "00101001" => data <= 768x"fffb87ffffd007ffffe007ff7f70177ffff00ffffff007fffff80ffff7f017fffff80ffffffc0ffffff80fff7f70077fffe007ffffc007ffffe803ffffd001f7ffd001ffffd001ffffc000ff7fd0017fffe000ffffc0007fffe000fffff0017f";
 when "00101010" => data <= 768x"fffb83fffff007ffffe007ff7f70077ffff807fffffc07fffffc0ffffffc17fffff80ffffffc07fffff807ff7f70077ffff003fffff401ffffe003ffff7011f7ffe001ffffc001ffffc000ff7fc0007fffe000fffff0007ffff000fffff0007f";
 when "00101011" => data <= 768x"fff883fffff007fffff803ff7f71077ffffc07fffffc07fffffc0ffffffc07fffffc0ffffffc07fffffc03ff7f7c07fffff803fffff001fffff001fffff011f7fff001fffff001ffffe000ff7f70007fffe000fffff0007ffff800fffff0007f";
 when "00101100" => data <= 768x"fffa83fffff001fffff803ff7f7c077ffffe03fffffc07fffffe0ffffff407fffffe07fffffc07fffffc03ff7f7c037ffff803fffffc01fffff803fffff011f7fff001fffff001ffffe000ff7ff0007fffe000fffff0007ffff800fffff0007f";
 when "00101101" => data <= 768x"fffffbfffffd41fffff803ff7f70037ffff807fffffc07fffffe0ffff7ff07fffffe0ffffffc07fffffc07ff7f7c077ffff803fffffc01fffff803fffff011f7ffe001fffff001ffffe000ff7f60017fffe000fffff000fffff800fff7f0047f";
 when "00101110" => data <= 768x"fffffffffff047fffff803ff7f70077ffff80ffffffc07fffffc0ffffff607fffffe0ffffffc07fffff807ff7f70077ffff803fffff017fffff003fffff01377ffe013ffffc011ffffe000ff7f4011ffffe001fffff001fffff008fffff005ff";
 when "00101111" => data <= 768x"fffbfffffff047fffff807ff7f70077ffff80ffffffc1ffffffc0ffffffc17fffffc0ffffffc07fffff80fff7f70077ffff007fffff007ffffe027fffff03777ffe023ffffc011ffffc003ff7fc011ffffe003ffffc011ffffe009ffff6005ff";
 when "00110000" => data <= 768x"fffbfffffff157fffff807ff7f71077ffff80ffffff41ffffff81ffffffc1ffffff81ffffff01ffffff80fff7f70077fffe007fffff047ffffe007ffffc047f7ffc027ffffc047ffffc003ff7fc0177fffc003ffffc017ffffc003ffffc013f7";
 when "00110001" => data <= 768x"fffffffffff1dffffff00fff7f70077ffff80ffffff01ffffff81ffffff01ffffff83ffffff41ffffff81fff7f701f7fffe00ffffff007ffffe007ffffc057f7ffc007ffffc047ffff8007ff7f40077fff8003ffffc007ffffc007ffffc017f7";
 when "00110010" => data <= 768x"fffffffffff1dffffff00fff7f70077ffff80ffffff01ffffff83ffffff03ffffff83ffffff01ffffff01fff7f701f7fffe00fffffc007ffffe00fffffc007f7ff8007ffffc007ffff8007ff7f00077fff8007ffffc007ffff800fffff8007f7";
 when "00110011" => data <= 768x"fffffffffff15fffffe00fff7f701f7ffff01ffffff01ffffff83ffffff07ffffff03ffffff07fffffe03fff7f701f7fffe01fffffc01fffffc00fffffc017f7ff800fffff0007ffff800fff7f00077fff800fffff001fffff800fffff001ff7";
 when "00110100" => data <= 768x"ffffffffffc55fffffe01fff7f701f7fffe03ffffff07ffffff03ffffff07ffffff03ffffff07fffffe03fff7f401f7fffe01fffffc01fffffc01fffffd01ff7ff800fffff000fffff800fff7f00177fff800fffff001fffff801fffff401ff7";
 when "00110101" => data <= 768x"ffffffffffc55fffffe01fff7f401f7fffe03fffffc07fffffe07ffff7f07ffffff07ffffff07fffffe03fff7f403f7fffe03fffffc01fffffc01fffffd01ff7ff800fffff000fffff800fff7f001f7fff800fffff001fffff801fffff401ff7";
 when "00110110" => data <= 768x"ffffffffffd55fffffe01fff7f401f7fffe03ffffff07fffffe07ffff7f07ffffff07ffffff07fffffe03fff7f701f7fffe03fffffc01fffffe01fffffc01ff7ff800fffff800fffff800fff7f001f7fff800fffff801fffffa00fffff401ff7";
 when "00110111" => data <= 768x"fffffffffff55fffffe00fff7ff01f7ffff03ffffff01ffffff03fffff707ffffff03ffffff01fffffe01fff7ff01f7fffe01fffffe41fffffe40fffffc417f7ffc007ffffc407ffff880fff7fc0077fff800fffffd007ffff800ffffff007f7";
 when "00111000" => data <= 768x"fffffffffff51fffffe00fff7f701f7ffff01ffffff01ffffff83ffffff07ffffff03ffffff01fffffe01fff7f701f7fffe00fffffc40fffffe00fffff5407f7ffe007ffffc407ffffc007ff7fc4077fffc807ffffd007ffffd007fffff007f7";
 when "00111001" => data <= 768x"fffffffffff75fffffe00fff7f701f7ffff01ffffff01ffffff81ffffff017fffff83ffffff01ffffff00fff7f70177fffe00fffffd007ffffe007ffffd007f7ffe203ffffc401ffffe003ff7f4403ffffe003ffffc407ffffe807fffff007f7";
 when "00111010" => data <= 768x"ffffffffffffdffffff80fff7f70177ffff00ffffffc1ffffff80ffffffc1ffffff81ffffffc1ffffff80fff7f7017fffff00ffffff007ffffe807fffff107ffffe003ffffc001ffffe003ff7f70017fffe003fffff401ffffe803fffff00777";
 when "00111011" => data <= 768x"fffffffffffdc7fffff00fff7ff0077ffff80ffffffc07fffffc0ffffffc1ffffffc0ffffffc0ffffff80fff7ff1077ffff007fffff007ffffe003fffff003ffffe003ffffc001ffffe001ff7ff001fffff001fffff401fffff801fffff001ff";
 when "00111100" => data <= 768x"fffffffffff547fffff807ff7f70077ffff80ffffffc07fffffc0ffffffc17fffffe0ffffffc07fffffc0fff7f7c077ffff803fffff017fffff003fffff011f7ffe001fffff001ffffe001ff7ff001fffff001fffff401fffff800fffff001ff";
 when "00111101" => data <= 768x"ffffe7fffffd47fffff807ff7f7c07fffffc07fffffc07fffffe0ffffffc17fffffe0ffffffc07fffffc07ff7f7c077ffff803fffff007fffff003ffff7011f7ffe001fffff001ffffe001ff7f7001fffff001fffffc01fffff800fffff001f7";
 when "00111110" => data <= 768x"fffffffffffdd7fffff803ff7f7c077ffffc07fffffc07fffffe0ffffff717fffffe0ffffffc07fffffe07ff7f7c077ffff803fffff007fffff003ffff7013f7ffe001ffffe001ffffe001ff7ff001fffff001fffff405fffff800fffff005f7";
 when "00111111" => data <= 768x"fffffffffffd57fffff807ff7ff0077ffff80ffffffc07fffffe0fffffff07fffffe0ffffffc07fffffc0fff7f74077ffff803fffff017fffff003fffff013f7ffe003ffffc001ffffe001ff7f7001fffff001fffff005fffff004fffff005f7";
 when "01000000" => data <= 768x"fffffffffff557fffff807ff7f7007fffff80ffffffc1ffffffc0ffffffc17fffffe0ffffffc1ffffff80fff7f70077ffff007fffff007ffffe027fffff007f7ffe023ffffc001ffffe003ff7f40117fffe003fffff001ffffe009fffff005f7";
 when "01000001" => data <= 768x"fffffffffff157fffff807ff7f7007fffff80ffffffc1ffffffc1ffffffc1ffffff81ffffffc1ffffff80fff7f70077ffff007fffff047ffffe007ffffd047f7ffe023ffffc047ffffc003ff7fc0177fffe003ffffc017ffffe00bffffc007f7";
 when "01000010" => data <= 768x"fffffffffff1fffffff00fff7f7007fffff80ffffff01ffffff81ffffff41ffffff81ffffffc1ffffff80fff7f701f7fffe00ffffff007ffffe007ffffc057f7ffc007ffffc047ffffc007ff7fc007ffffc007ffffc017ffffc007ffffc017f7";
 when "01000011" => data <= 768x"fffffffffff5fffffff00fff7f7007fffff00ffffff01ffffff81ffffff01ffffff83ffffff01ffffff01fff7f701f7fffe00fffffe007ffffe00fffffc007f7ffc007ffffc047ffff8007ff7fc0077fff8007ffffc007ffff800fffffc017f7";
 when "01000100" => data <= 768x"fffffffffff15ffffff007ff7f7007fffff80ffffff01ffffff81ffffff01ffffff81ffffff81ffffff81fff7f701f7ffff00ffffff007ffffe007fff7f007f7ffe003ffffc007ffff8003ff7f40037fff8003ffffc007ffff8007ffffc007f7";
 when "01000101" => data <= 768x"fff3fffffff047fffff003ff7f70077ffff807fffff007fffff80ffffffc1ffffff80ffffffc1ffffff80fff7f70077ffff007fffff007ffffe003fff7f013ffffe003ffffc011ffffc001ff7fc011ffff8000ffffc001ffffc000ffffc001ff";
 when "01000110" => data <= 768x"fff0fffffff041fffff001ff7f7001fffff803fffff005fffff803fffffc07fffff807fffffc07fffff807ff7f70077ffff803fffff005ffffe001fff7f001fffff000fffff0047fffe0087f7f70047fffe0003fffc0041fffc0003fffc0041f";
 when "01000111" => data <= 768x"fffbfffffff050fffff000ff7f70007ffff800fffffc01fffff803fffffc01fffff803fffffc03fffff803ff7f7407fffff803fffff401fffff801fffff0017ffff0007ffff0007ffff8003f7f70041ffff8021ffff0071fffe0020fff70031f";
 when "01001000" => data <= 768x"fffa383ffff0007ffff8003f7f7c003ffff8003ffffc007ffffc007ffffc007ffffc00fffffc01fffff800ff7f7d01fffffa01fffffc01fffffc00fffffc007ffffe003ffffc001ffffc000f7f740117fffe0307fffc0107fff80103fff00103";
 when "01001001" => data <= 768x"ffff0a1ffffc001ffffe000f7f7f011ffffe000ffffc001ffffe001fffff0017ffff000fffff001ffffe803f7f7f007ffffe003fffff007ffffe007ff7f7007fffff003fffff0017fffe00077f770007fffe0003ffff0101fffe0081fffc0111";
 when "01001010" => data <= 768x"fffffe1fffffc01fffff800f7f7f0007ffff000fffff000fffff000ff7f70007ffff8007ffffc007ffff800f7f7f9007ffff800fffffc00fffff800ff7ff801fffff803fffff001fffff000f7f7f0017ffff0003ffff0005ff9e0001f7000041";
 when "01001011" => data <= 768x"fffffe3ffffff41fffffe03f7f7fc01fffff800fffff000fffff800fffff0007ffff8007ffffc007ffffc0077f7f4007ffffe007ffffc007ffffe007fff7c017ffffc00fffffc01fffff801f7f5f0017ff0f8007ff040007ff000007ff000007";
 when "01001100" => data <= 768x"fffffffffffffc7ffffff8ff7f7f711fffffc01fffffc01fffff800fffff0017ffff800fffffc007ffffc0077f7f4007ffffe007fffff007ffffe007fff7f017ffffe00fffdfc05fff8f803f7f074037ff80002fffc0001fffe0000ffff00017";
 when "01001101" => data <= 768x"fffffffffffff1fffffff8ff7f7f707fffffc03fffffc01fffff801fffff001fffff800fffffc01fffffc00f7f7f4007ffffe00ffffff007ffffe00ffffff017ffefe03fff07c05fff87c03f7f01003fff80002ffff0001ffff0001ffff0001f";
 when "01001110" => data <= 768x"fffffffffffff1fffffff1ff7f7f717fffffc03fffffc01fffff801fffff001fffff800fffffc01fffffc00f7f7f401fffffe00ffffff01fffffe00fffd7f01fff8fe03fff07c07fff83803f7f41003fffe0003ffff0001fffe0001ffff0001f";
 when "01001111" => data <= 768x"fffffffffffff7ffffffe3ff7f7f717fffffc03fffff801fffff803fffff001fffff001fffffc01fffffc01f7f7fc01fffffe01fffffe01fffffe01fffd7f01fff8fe03fff07c07fff80803f7fd0003fffe0001fffe0001fffe0003fffc0001f";
 when "01010000" => data <= 768x"fffffffffffff7ffffffe3ff7f7f717fffff803fffff005fffff003fffff001fffff001fffff401fffff801f7f7fc01fffffe01fffffc01fffffe01fff57f05fff8f803fff05c07fff80803f7fd0007fffe0003fffc0001fffe0003fffc0001f";
 when "01010001" => data <= 768x"ffffffffffffd7ffffffe7ff7f7fc07fffff807fffff007fffff003fffff0017ffff003fffff001fffff801f7f7fc01fffffe03fffffc01fffffe01fff57f05fff8f807fff05c07fff80807f7fd0007fffe0003fffc0001fffe0003fffc0001f";
 when "01010010" => data <= 768x"ffffffffffffffffffffc7ff7f7f417fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff8f807fff05c07fff80807f7fd0007fffe0003fffc0005fffe0003fffc0001f";
 when "01010011" => data <= 768x"ffffffffffffffffffffc7ff7f7f417fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff8f807fff07c07fff80807f7fd0007fffe0003ffff0005fffe0003fffe00017";
 when "01010100" => data <= 768x"ffffffffffffd7ffffffc7ff7f7fc07fffff807fffff007fffff003fffff0037ffff003fffff001fffff803f7f7fc01fffffc03fffffc01fffffe03fff57e05fff87a07fff05c07fff80807f7fd0007fffe0003ffff0005fffe0003ffff00017";
 when "01010101" => data <= 768x"ffffffffffffd7ffffffc3ff7f7fc07fffff807fffff007fffff003fffff0017ffff003fffff001fffff801f7f7fc01fffffc01fffffc01fffffe03fff47e07fff87e07fffc5c07fff80807f7fd0007fffe0003ffff0005fffe0003ffff00017";
 when "01010110" => data <= 768x"ffffffffffffc7ffffffc2ff7f7fc07fffff803fffff007fffff003fffff001fffff003fffff001fffff801f7f7fc01fffffc01fffffc01fffefe01fffc7e05fff87e03fffc5c07fffc0807f7ff0007ffff0003ffff0005fffe0003ffff00017";
 when "01010111" => data <= 768x"ffffffffffffc7ffffffc0ff7f7fc07fffff803fffff005fffff003fffff001fffff001fffff001fffff801f7f7fc01fffffc01fffffc01fffefe00fffc7e01fff83e03fffc5c07fffc0807f7ff0007ffff0003ffff0005fffe0003ffff00017";
 when "01011000" => data <= 768x"ffffefffffffc7ffffffe0ff7f7fc07fffff803fffff001ffffe001fffff001fffff001fffff001fffff800f7f7fc01fffffc00fffffc01fffe7e00fffc7e01fff83e03fffc1c07fffe0803f7f70007ffff0003ffff0001fffe0001ffff0001f";
 when "01011001" => data <= 768x"ffffe7ffffffc5ffffffe07f7f7fc07fffff803fffff001ffffe001fffff001fffff000fffff001fffff800f7f7fc017ffffc00fffffc01fffe3e00fffc1e017ffc3e03fffc1c05fffe0803f7f70003ffff0003ffff00017ffe0000ffff0001f";
 when "01011010" => data <= 768x"ffffe3ffffffc17fffffe03f7f7f401fffff003fffff001ffffe001fffff001fffff000fffff000fffff800f7f7f4007ffffc00ffff7c007ffe3e00fffc1e017ffc3e03fffc1c05fffe0803f7f70003ffff0003ffff00017ffe0000ffff0001f";
 when "01011011" => data <= 768x"ffffe3ffffffc17fffffe03f7f7f401fffff001fffff001ffffe000fffff0017ffff000fffff0007ffff800f7fff4007ffffc00ffff5c007ffe1e00fffc1e017ffe1e01fffc0401ffff0003f7f70001ffff0003ffff00017fff0000ffff00017";
 when "01011100" => data <= 768x"ffffe1fffffff17fffffe03f7f7f001fffff001fffff001ffffe000fffff0007ffff0007ffff0007ffff80077fff4007ffffc007fff5c007ffe0e007ffc1e017ffe0e01ffff0401ffff8003f7f70001ffff0001ffff0001ffff00003fff01017";
 when "01011101" => data <= 768x"ffffe1fffffff05fffffc01f7f7f001fffff000fffff0007fffe000fffff0007ffff0007ffff4007ffff80077fffc007ffffc007fff1c007ffe0e007fff17017ffe0e00ffff0401ffff8003f7ff0001ffff8001ffff0001ffff0000bfff01007";
 when "01011110" => data <= 768x"ffffe0fffffff01fffffc01f7f7f001fffff000fffff0007fffe0007ffff0007ffff0007ffff4007ffff80077f7fc007fffbc003fff0c007ffe0e003fff07017fff0600bfff0401ffff8000f7ff0001ffff8001ffff0001ffff8000bfff01007";
 when "01011111" => data <= 768x"fffff0fffffff01fffffc00f7f7f001fffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7fc007fffac003fff04007ffe0e003fff07017fff0200bfff44017fff8000f7f740017fff8001ffff0001ffff8000bfff00017";
 when "01100000" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0017ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7fc007fff8c003fff04007fff06003fff07003fff0200bfffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "01100001" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0017ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "01100010" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007ffff0007ffff0003ffff4007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "01100011" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007ffff0007ffff0003ffff0007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff04011";
 when "01100100" => data <= 768x"fffff0ffffffd01fffffc00f7f7f0007ffff000fffff0007fffe0007fff70007ffff0003ffff0007ffff80037f7f4007fff84003fff04007fff06003fff07003fff82003fffc0005fffc000f7f7c0017fff8001ffffc001ffff8000ffff05011";
 when "01100101" => data <= 768x"fffff0ffffffd05fffffc00f7f7f001fffff000fffff0007fffe0007fff70007ffff0003ffff0007ffff80037f7f0007fff84003fff04007fff06003fff06003fff82003fffc0007fffc000f7f7c0017fff8001ffff0001ffff8000ffff04011";
 when "01100110" => data <= 768x"fffff0fffffff05fffff800f7f7f001fffff000fffff0007fffe0007ffff0007ffff0003ffff0007ffff80037f7f0007fff88003fff04007fff06003fff06003fff02003fffc0007fff8000f7ff40017fff8001ffff0001ffff8000ffff04011";
 when "01100111" => data <= 768x"fffff0fffffff05fffff800f7f7f001fffff000fffff0007fffe0007ffff0007fffe0007ffff0007ffff80037f7f0007fff8c003fff04007ffe06003fff04003fff0200bfff40007fff8000f7f780017fff8001ffff0001ffff8000ff7f04011";
 when "01101000" => data <= 768x"ffffe0ffffffd05fffff801f7f7f001ffffe000fffff0007fffe000ffffc0007fffe0007ffff0007ffff80037f7f0007fff88003fff04007ffe0e003fff04017fff0600bfff04007fff8000f7f710017fff8001ffff0001ffff8000ffff04011";
 when "01101001" => data <= 768x"ffffe0ffffffd05fffff801f7f7f001ffffe000ffffc0007fffe000ffffc0007fffe0007ffff0007ffff80077f7f0007fffb8003fff04007ffe0c003fff04017fff0600bfff04017fff8000f7f71001ffff8001ffff0001ffff8000ffff04001";
 when "01101010" => data <= 768x"ffffc3ffffffc07fffff803f7f7f011ffffe001ffffc001ffffc000ffffc0007fffe0007fffd0007ffff00077f7f0007fffb8007fff1c007ffe0c007fff14017ffe0e00bfff0401ffff8000f7ff1001ffff0001ffff0001ffff0000ffff04011";
 when "01101011" => data <= 768x"ffff83ffffffc07fffff803f7f7f011ffffe001ffffc001ffffc000ffffc0017fffc000ffffc0007ffff000f7fff0007ffff8007ffd1c007ffe0c007ffc1c017ffe0c00ffff0401ffff8000f7ff0001ffff0001ffff0001ffff0000ffff10011";
 when "01101100" => data <= 768x"ffff03ffffff807fffff803f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc000fffff000f7f7f0007ffff000fffd5d007ffe1800fffc1d017ffe0c03fffc0401fffe0001f7f70001ffff0003ffff0001ffff0001fff700017";
 when "01101101" => data <= 768x"ffff02ffffff007fffff803f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc001ffffe000f7fff0017ffff800ffff7901fffe3900fffc11017ff81a03fffc1c01fffc0801f7f70001ffff0003ffff0001fffe0001ffff00017";
 when "01101110" => data <= 768x"fffe00ffffff007fffff003f7f7f003ffffe003ffffc001ffffc001ffffc001ffff8000ffffc001ffffe000f7fff001fffff800fffff901fffff980fffd71017ff83a03fffc1c01fff81801f7fc0001fffe0003ffff0001ffff0003ffff00017";
 when "01101111" => data <= 768x"fff800fffffc007ffffe007f7f7c003ffffc003ffffc001ffff8001ffff8001ffff8000ffffc001ffffe000f7f7f001fffff800fffff101fffff880ffff71017ffaf803fff07c01fff07803f7f07c01fff80803fffc0001fffe0003fff700017";
 when "01110000" => data <= 768x"ffe001fffff001fffff000ff7ffd007ffff8003ffff0001ffff8003ffff0001ffff0001ffff0001ffff8000f7f7f001fffff001fffff005fffff800fffff1037ffffa03fffffc01fffff800f7f1fc11ffe1f800ffc1fc01ffc0a800ff400001f";
 when "01110001" => data <= 768x"ffe303ffffc001ffffc000ff7f70017ffff0007ffff0007ffff0003ffff0001ffff0003ffff0001ffff0001f7f75001fffff001fffff101ffffe000ffff7501fffff201fffff401fffff800f7f7f4017ffffc007ffffc017ffbfc003fc17c013";
 when "01110010" => data <= 768x"ffffe7ffffd541ffffc001ff7fc0017fffe0007ffff0007ffff8003ffff0013ffff0003ffff0001ffff0001f7f70001ffffa001fffff001ffffe000fffff501ffffe581ffffc501ffffee00f7f7f4007ffffe007ffff4007ffffe003ffffc001";
 when "01110011" => data <= 768x"fffffffffffffdfffffee0ff7f70007ffff0003ffff0005ffffc003ffffc001ffff8001ffffc001ffff8000f7f7c001ffff8000ffffd000fffff000fffff4017fffe080fffff5c07fffe78077f7f5007fffef803fffff001fffff001fffff001";
 when "01110100" => data <= 768x"ffffffffffffffffffffffff7f7fc51fffff800fffffc007ffff800fffff0007ffff0007ffff0007fffe00037f7f0007ffff0003ffff4007ffffc003fff7c007ffffc003ffffc407ffff8e037f7f1f01ffffbe00ffff7c00fffffc00fffffc00";
 when "01110101" => data <= 768x"fffffffffffffffffffffe3f7f7f7f17fffffe03fffff401fffff000fffff001ffffe000ffffc000ffffc0007f7fc000fffff000fffff000fffff000fffff000fffff800fffff100fffffb007f7f7701fffff700ffffff00ffffff00fffff700";
 when "01110110" => data <= 768x"fffffff0fffffff0ffffff807f7f7f00fffffe00fffffc00fffffc00fffffc00fffffc00fffffc00fffffe007f7f7700fffffe00ffffff00fffffe00ffffff40ffffff80ffffffc0ffffff807f7f7fc0ffffff80ffffffc0ffffff80fffff790";
 when "01110111" => data <= 768x"fffffffffffffff4ffffffe07f7f7f41ffffff80ffffffc0ffffff80ffffffc0ffffffc0ffffffc0ffffffc07f7f7f40ffffffe0ffffffd0ffffffc0ffffff40ffffffc0ffffffc0ffffffc07f7f7f00ffffff00fffffd00fffffe00fffff400";
 when "01111000" => data <= 768x"fffffffffffffffdfffffff87f7f7f71fffffff0fffffff0fffffff0f7f7fff0fffffff0fffffff0fffffff0757f7f74fa3ffff8f4557c40f0202800f0400000f0200000f5400100ffe002007f500700ffe00200ffc00100ffe00000ffd00100";
 when "01111001" => data <= 768x"ffff0fffffff57ffffff8fff777f477ffeba03fff50007fffe0003fefd0001f5ff0003f8ff0001f4ff8000f87f400170ff800020ffc00000ffe00000f7701510fff03f80fff47dc0ffffff807f777f00ffffff00ffffff00ffffff00f7f7f700";
 when "01111010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f5fffffffbffffffd5ffffffbaffffff557fffff23fffffd55fffffe03f7f7f517fffff803fffff407fffff803fffff0037";
 when "01111011" => data <= 768x"fffbffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01111100" => data <= 768x"fff03ffffff07ffffff8ffff7f7d7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01111101" => data <= 768x"fffffffffff07ffffff03fff7ff11f7ffff03ffffff01ffffffc7fffffff7fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01111110" => data <= 768x"ffffffffffffffffffffffff7f7d7f7ffff81ffffff01ffffff80ffffff01ffffff81ffffffc7fffffffffff7f7fff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "01111111" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffff5ffffffc1ffffff41ffffff80ffffff00ffffff80fff7f7c1f7ffffe3fffffff7fffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10000000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff7ffffffe3ffffffc1ffffffc0fff7f7c077ffff807fffffc07fffffc0fffffff5fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10000001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffffffffffffffffffffffffffe0fff7f7c077ffff807fffffc07fffff807fffff407fffffe0fffffff5fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10000010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f5f7ffffe0ffffffc07fffffc07fffffc07fffff803fffffc07fffffe0fff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10000011" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7fffffbfffffff1ffffffc07fffffc07fffff803fffffc07fffffc07ff7f7c07ffffff3ffffffffffffffffffffffff7ff";
 when "10000100" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7fff7fffffffffffff17fffffc07fffffc07fffff803fffffc05fffffc07ff7f7c077fffff0fffffffdfffffffffffffffffff";
 when "10000101" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f7f7fffff3ffffffc07fffffc07fffffc07fffff803fffffc07fffffc07ff7f7f177fffff3ffffffffffffffffffffffff7ff";
 when "10000110" => data <= 768x"ffffffffffffffffffffffff7fff7f7fffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f177ffffe07fffffc07fffff803fffffc07fffff803fffffc07fffffe0fff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10000111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffffffffffff1ffffffe0fff7f74077ffff803fffffc07fffff803fffffc07fffffe0fffffff5fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff7ffffffe0ffffffc07fffff807ff7f70077ffff803fffff407fffffc0ffffff51fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffe3ffffffc17fffff807fffff007fffff807ff7f7107fffff807fffffc07fffffe9fffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001010" => data <= 768x"ffffffffffffffffffffffff7f7fff7ffffffffffffd5ffffffc0ffffff017fffff007fffff007fffff807ff7f70077ffff80ffffffc5ffffffeefffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001011" => data <= 768x"ffffffffffffffffffffffff7f7fff7fffffffffffff5ffffffc0ffffff007fffff807fffff007fffff003ff7f70077ffff80ffffffc1fffffffbffffff7ffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001100" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffff7ffffffe1ffffffc07fffff807fffff007fffff803ff7f7003fffff807fffffc07fffffe3fffffffffffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001101" => data <= 768x"ffffffffffffffffffffffff7f7fff7fffffffffffffdfffffffbffffffc17fffff803fffff801fffff803ff7f7803fffff803fffffc07fffffe0fffffff5fffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001110" => data <= 768x"ffffffffffffffffffffffff7f7fff7ffffffffffffffffffffffffffffd07fffffe03fffffc01fffff803ff7f71017ffff803fffffc01fffffe07ffffff17ffffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10001111" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffff57fffffe03fffffc01fffffc01ff7f7c01fffff801fffffc01fffffc03fffff407ffffff2fffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010000" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffffff7ffffff83fffffd05fffffc01ff7f7c01fffff801fffffc01fffffc01fffff401ffffff03ffffff57ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010001" => data <= 768x"ffffffffffffffffffffffff7f7f7f7ffffffffffffffffffffffffffff7ffffffffafffffff05fffffe01ff7f7c01fffffc01fffffc01fffffc01fffff401fffffe03ffffff57ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010010" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffbfffffff07fffffc03ff7f7c017ffff801fffffc01fffffc01fffff407fffffe03ffffff1dffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010011" => data <= 768x"ffffffffffffffffffffffff7f7f7f7fffffffffffffffffffffffffffffffffffffffffffff07fffffc03ff7f7c017ffff803fffffc01fffff803fffffc117ffffe03ffffff47ffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010100" => data <= 768x"ffa00000fffd5555ffffffff7f7ffffffffffffffffffffffffffffffff7fff7fffffffffffc07fffffc03ff7f7c037ffff803fffffc01fffff803fffffc07f7fffc07fffffd1fffffffffff7f7f7f7fffffffffffffffffffffffffffffffff";
 when "10010101" => data <= 768x"20000000d5540000fffc00007f7c0001fffe0000ffff5400fffffe00f7ffff11fffffe03ffff0505fffc06037f740701fff80380fff40741fff80380f7fc0751fffc07f2fffd1fd5fffffffa7f7f7f77ffffffffffffffffffffffffffffffff";
 when "10010110" => data <= 768x"022bffff0005ffff0007ffff0007ff7f0003ffff0001c17f0000e07f0001c0770001e03e0001f01c0003f80800077800000ff8000007fc000007fc000007fc000003f8000001f000000020000000000000000000000000000000000000000000";
when others => data <= 768x"0";
end case;
end if;
end process;
end;
